netcdf leorgn_ysi_blue_green_algae {
dimensions:
	feature_type_instance = 1 ;
	time = UNLIMITED ; // (4040 currently)
	height = 1 ;
	text = 128 ;
variables:
	char platform(text) ;
		platform:imo_code = "" ;
		platform:ioos_code = "urn:ioos:station:glos:leorgn" ;
		platform:call_sign = "" ;
		platform:ices_code = "" ;
		platform:long_name = "Oregon Pump Station" ;
        platform:wmo_code = "" ;
		platform:short_name = "Oregon_Pump_Station" ;
	int crs ;
		crs:inverse_flattening = 298.257223563 ;
		crs:epsg_code = "EPSG:4326" ;
		crs:long_name = "http://www.opengis.net/def/crs/EPSG/0/4326" ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:semi_major_axis = 6378137. ;
	char feature_type_instance(text) ;
		feature_type_instance:cf_role = "timeseries_id" ;
		feature_type_instance:long_name = "Identifier for each feature type instance" ;
	double time(time) ;
		time:time_coverage_end = "2017-08-31T23:50:00+0000" ;
		time:time_coverage_start = "2017-08-01T00:00:00+0000" ;
		time:calendar = "gregorian" ;
		time:units = "seconds since 1970-01-01T00:00:00Z" ;
		time:standard_name = "time" ;
		time:long_name = "time of measurement" ;
		time:axis = "T" ;
	char instrument(text) ;
		instrument:serial_number = "" ;
		instrument:comment = "" ;
		instrument:calibration_date = "" ;
		instrument:definition = "http://mmisw.org/ont/ioos/definition/sensorID" ;
		instrument:long_name = "urn:ioos:sensor:glos:leorgn:ysi_blue_green_algae" ;
		instrument:make_model = "" ;
	double longitude ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "sensor longitude" ;
		longitude:axis = "X" ;
	double latitude ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "sensor latitude" ;
		latitude:axis = "Y" ;
	double obs(time, feature_type_instance) ;
		obs:instrument = "instrument" ;
		obs:nc_name = "leorgn_ysi_blue_green_algae.nc" ;
		obs:scale_factor = 1. ;
		obs:short_name = "YSI Blue Green Algae" ;
		obs:nodc_name = "" ;
		obs:_FillValue = -9999. ;
		obs:target = "/tmp/leorgn_ysi_blue_green_algae" ;
		obs:add_offset = 0. ;
		obs:platform = "platform" ;
		obs:habs_name = "blue_green_algae" ;
        obs:long_name = "ysi_blue_green_algae" ;
		obs:standard_name = "blue_green_algae" ;
		obs:featureType = "timeSeries" ;
		obs:units = "1" ;
		obs:keywords = "EARTH SCIENCE > BIOLOGICAL CLASSIFICATION > PLANTS > MICROALGA" ;
		obs:depth = 0. ;
		obs:source = "platform/leorgn/leorgn_ysi_blue_green_algae" ;
		obs:keywords_vocabulary = "GCMD Earth Science Keywords. Version 5.3.3" ;
		obs:coverage_content_type = "physicalMeasurement" ;
		obs:grid_mapping = "crs" ;
		obs:coordinates = "time latitude longitude height" ;
	double height(height) ;
		height:positive = "down" ;
		height:units = "m" ;
		height:long_name = "height of the sensor relative to sea surface" ;
		height:standard_name = "height" ;
		height:axis = "Z" ;

// global attributes:
        :contributor_name = "GLOS" ;
        :contributor_role = "Data Provider" ;
        :creator_country = "USA" ;
        :creator_email = "example@gmail.com" ;
		:creator_sector = "academic" ;
        :instrument = "instrument" ;
        :comment = "test data" ;
        :geospatial_vertical_units = "" ;
        :geospatial_lat_max = 41.67196 ;
        :Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
        :project = "" ;
        :creator_name = "Bob" ;
        :creator_phone = "401 783 9999" ;
        :geospatial_vertical_resolution = "" ;
        :time_coverage_end = "" ;
        :time_coverage_duration = "" ;
        :date_modified = "201791" ;
        :geospatial_lat_units = "degrees_north" ;
        :nodc_template_version = "NODC_NetCDF_TimeSeries_Orthogonal_Template_v1.1" ;
        :featureType = "timeSeries" ;
        :publisher_name = "GLOS" ;
        :date_created = "201791" ;
        :time_coverage_resolution = "" ;
        :title = "Oregon Pump Station" ;
        :cdm_data_type = "station" ;
        :geospatial_lon_resolution = "" ;
        :acknowledgment = "" ;
        :geospatial_vertical_min = "" ;
        :standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention Standard Name Table v26" ;
        :publisher_email = "dmac@glos.us" ;
        :missing_value = -9999. ;
        :source = "" ;
        :references = "" ;
        :geospatial_lon_max = -83.2903 ;
        :Conventions = "CF-1.6" ;
        :geospatial_lat_resolution = "" ;
        :history = "" ;
        :metadata_link = "" ;
        :creator_url = "www.example.com" ;
        :creator_address = "123 Main St" ;
        :creator_city = "Lansing" ;
        :creator_state = "Michigan" ;
        :creator_zipcode = "01532" ;
        :naming_authority = "GLOS" ;
        :date_issued = "201791" ;
        :geospatial_lon_min = -83.2903 ;
        :license = "Freely Distributed" ;
        :institution_dods_url = "" ;
        :geospatial_vertical_max = "" ;
        :time_coverage_start = "" ;
        :uuid = "" ;
        :keywords_vocabulary = "" ;
        :institution_url = "http://glos.us" ;
        :id = "leorgn" ;
        :keywords = "EARTH SCIENCE > BIOLOGICAL CLASSIFICATION > PLANTS > MICROALGA" ;
        :platform = "platform" ;
        :geospatial_lon_units = "degrees_east" ;
        :sea_name = "Great Lakes" ;
        :institution = "GLOS, City of Oregon, Ohio, Oregon Pump Station" ;
        :geospatial_vertical_positive = "" ;
        :summary = "Data from Great Lakes Oregon Pump Station" ;
        :publisher_url = "http://glos.us" ;
        :publisher_country = "USA" ;
        :publisher_address = "123 Main St." ;
        :publisher_city = "Lansing" ;
        :publisher_state = "Michigan" ;
        :publisher_zipcode = "01532" ;
        :publisher_phone = "401 783 9999" ;
		:geospatial_lat_min = 41.67196 ;
		:processing_level = "none" ;
        :platform_vocabulary = "https://mmisw.org/orr/#http://mmisw.org/ont/ioos/platform" ;
}
