netcdf ooi_glider {
dimensions:
    obs = 2;
    maxStrlen64 = 64 ;
    traj = 1 ;
variables:
    char trajectoryId(traj, maxStrlen64) ;
        trajectoryId:long_name = "trajectory identifier" ;
        trajectoryId:cf_role = "trajectory_id" ;
    int nobs(traj) ;
        nobs:long_name = "number of obs for this profile" ;
        nobs:sample_dimension = "obs" ;
    double time(obs) ;
        time:units = "seconds since 1900-01-01 0:0:0" ;
        time:long_name = "time of measurement" ;
    double latitude(obs) ;
        latitude:units = "degrees_north" ;
        latitude:long_name = "latitude of measurement" ;
    double longitude(obs) ;
        longitude:units = "degrees_east" ;
        longitude:long_name = "longitude of measurement" ;
    double altitude(obs) ;
        altitude:units = "m" ;
        altitude:long_name = "altitude of measurement" ;
        altitude:positive = "up" ;
    float m_present_secs_into_mission(obs) ;
        m_present_secs_into_mission:units = "s" ;
        m_present_secs_into_mission:long_name = "Elapsed mission time, Secs" ;
        m_present_secs_into_mission:_FillValue = -9999999.f ;
        m_present_secs_into_mission:comment = "Secs since mission started" ;
        m_present_secs_into_mission:coordinates = "time latitude longitude altitude" ;
    double ingestion_timestamp(obs) ;
        ingestion_timestamp:units = "seconds since 1900-01-01" ;
        ingestion_timestamp:long_name = "Ingestion Timestamp, UTC" ;
        ingestion_timestamp:coordinates = "time latitude longitude altitude" ;
        ingestion_timestamp:_FillValue = -9999. ;
        ingestion_timestamp:comment = "The NTP Timestamp for when the granule was ingested" ;
    double port_timestamp(obs) ;
        port_timestamp:units = "seconds since 1900-01-01" ;
        port_timestamp:long_name = "Port Timestamp, UTC" ;
        port_timestamp:_FillValue = -9999999. ;
        port_timestamp:comment = "Port timestamp, UTC" ;
        port_timestamp:coordinates = "time latitude longitude altitude" ;
    double sci_seawater_density(obs) ;
        sci_seawater_density:units = "kg m-3" ;
        sci_seawater_density:long_name = "Seawater Density" ;
        sci_seawater_density:coordinates = "time latitude longitude altitude" ;
        sci_seawater_density:data_product_identifier = "DENSITY_L2" ;
        sci_seawater_density:standard_name = "sea_water_density" ;
        sci_seawater_density:_FillValue = -9999999. ;
        sci_seawater_density:comment = "The density of seawater in kg m-3 computed using the TEOS-10 equations with data from the conductivity, temperature and depth (CTD) family of instruments." ;
    float sci_water_pressure(obs) ;
        sci_water_pressure:units = "bar" ;
        sci_water_pressure:long_name = "Seawater Pressure" ;
        sci_water_pressure:_FillValue = -9999999.f ;
        sci_water_pressure:comment = "Seawater Pressure refers to the pressure exerted on a sensor in situ by the weight of the column of seawater above it. It is calculated by subtracting one standard atmosphere from the absolute pressure at the sensor to remove the weight of the atmosphere on top of the water column. The pressure at a sensor in situ provides a metric of the depth of that sensor. Units: bar" ;
        sci_water_pressure:coordinates = "time latitude longitude altitude" ;
    float sci_m_present_secs_into_mission(obs) ;
        sci_m_present_secs_into_mission:units = "s" ;
        sci_m_present_secs_into_mission:long_name = "Elapsed mission time based on science derived start time, Secs" ;
        sci_m_present_secs_into_mission:_FillValue = -9999999.f ;
        sci_m_present_secs_into_mission:comment = "Secs since mission started. Based on Science derived start time." ;
        sci_m_present_secs_into_mission:coordinates = "time latitude longitude altitude" ;
    double sci_water_pracsal(obs) ;
        sci_water_pracsal:units = "1" ;
        sci_water_pracsal:long_name = "Practical Salinity" ;
        sci_water_pracsal:_FillValue = -9999999. ;
        sci_water_pracsal:comment = "Salinity is generally defined as the concentration of dissolved salt in a parcel of seawater. Practical Salinity is a more specific unitless quantity calculated from the conductivity of seawater and adjusted for temperature and pressure. It is approximately equivalent to Absolute Salinity (the mass fraction of dissolved salt in seawater) but they are not interchangeable. Units: unitless" ;
        sci_water_pracsal:data_product_identifier = "PRACSAL_L2" ;
        sci_water_pracsal:standard_name = "sea_water_practical_salinity" ;
        sci_water_pracsal:coordinates = "time latitude longitude altitude" ;
    char preferred_timestamp(obs, maxStrlen64) ;
        preferred_timestamp:units = "1" ;
        preferred_timestamp:long_name = "Preferred Timestamp" ;
        preferred_timestamp:_FillValue = "e" ;
        preferred_timestamp:comment = "Timestamp preferred as official record." ;
        preferred_timestamp:coordinates = "time latitude longitude altitude" ;
    double sci_ctd41cp_timestamp(obs) ;
        sci_ctd41cp_timestamp:units = "seconds since 1970-01-01" ;
        sci_ctd41cp_timestamp:long_name = "Ctd41cp Timestamp, UTC" ;
        sci_ctd41cp_timestamp:_FillValue = -9999999. ;
        sci_ctd41cp_timestamp:comment = "CTD41CP Timestamp in seconds since January 01, 1970. UTC" ;
        sci_ctd41cp_timestamp:coordinates = "time latitude longitude altitude" ;
    char provenance(obs, maxStrlen64) ;
        provenance:name = "provenance" ;
        provenance:coordinates = "time latitude longitude altitude" ;
    float sci_water_temp(obs) ;
        sci_water_temp:units = "deg_C" ;
        sci_water_temp:long_name = "Seawater Temperature" ;
        sci_water_temp:data_product_identifier = "TEMPWAT_L1" ;
        sci_water_temp:standard_name = "sea_water_temperature" ;
        sci_water_temp:coordinates = "time latitude longitude altitude" ;
        sci_water_temp:_FillValue = -9999999.f ;
        sci_water_temp:comment = "Seawater temperature near the sensor. Units: degrees Celsius" ;
    double internal_timestamp(obs) ;
        internal_timestamp:units = "seconds since 1900-01-01" ;
        internal_timestamp:long_name = "Internal Timestamp, UTC" ;
        internal_timestamp:coordinates = "time latitude longitude altitude" ;
        internal_timestamp:_FillValue = -9999999. ;
        internal_timestamp:comment = "Internal timestamp, UTC" ;
    char quality_flag(obs, maxStrlen64) ;
        quality_flag:name = "quality_flag" ;
        quality_flag:coordinates = "time latitude longitude altitude" ;
    float sci_water_cond(obs) ;
        sci_water_cond:units = "S m-1" ;
        sci_water_cond:long_name = "Seawater Conductivity" ;
        sci_water_cond:_FillValue = -9999999.f ;
        sci_water_cond:comment = "Seawater conductivity refers to the ability of seawater to conduct electricity. The presence of ions in the seawater, such as salt, increases the electrical conducting ability of seawater. As such, conductivity can be used as a proxy for determining the quantity of salt in a sample of seawater. Units: S m-1" ;
        sci_water_cond:coordinates = "time latitude longitude altitude" ;
        sci_water_cond:data_product_identifier = "CONDWAT_L1" ;
        sci_water_cond:standard_name = "sea_water_electrical_conductivity" ;
    double driver_timestamp(obs) ;
        driver_timestamp:units = "seconds since 1900-01-01" ;
        driver_timestamp:long_name = "Driver Timestamp, UTC" ;
        driver_timestamp:_FillValue = -9999999. ;
        driver_timestamp:comment = "Driver timestamp, UTC" ;
        driver_timestamp:coordinates = "time latitude longitude altitude" ;
    char id(obs, maxStrlen64) ;
        id:name = "id" ;
        id:coordinates = "time latitude longitude altitude" ;
    double m_present_time(obs) ;
        m_present_time:units = "seconds since 1970-01-01" ;
        m_present_time:long_name = "Time at the start of the cycle, UTC" ;
        m_present_time:_FillValue = -9999999. ;
        m_present_time:comment = "Secs since 1970 @ start of cycle" ;
        m_present_time:coordinates = "time latitude longitude altitude" ;
    int deployment(obs) ;
        deployment:name = "deployment" ;
        deployment:coordinates = "time latitude longitude altitude" ;
    double sci_m_present_time(obs) ;
        sci_m_present_time:units = "seconds since 1970-01-01" ;
        sci_m_present_time:long_name = "Science derived time at the start of the cycle, UTC" ;
        sci_m_present_time:coordinates = "time latitude longitude altitude" ;
        sci_m_present_time:_FillValue = -9999999. ;
        sci_m_present_time:comment = "Written by science on every cycle their notion of time, secs since 1970" ;

// global attributes:
        :Conventions = "CF-1.6" ;
        :history = "2016-06-14T16:07:44.373980 generated from Stream Engine" ;
        :node = "GL340" ;
        :comment = "" ;
        :publisher_email = "" ;
        :sourceUrl = "http://oceanobservatories.org/" ;
        :collection_method = "telemetered" ;
        :stream = "ctdgv_m_glider_instrument" ;
        :featureType = "trajectory" ;
        :creator_email = "" ;
        :publisher_name = "Ocean Observatories Initiative" ;
        :date_modified = "2016-06-14T16:07:44.374181" ;
        :keywords = "" ;
        :cdm_data_type = "trajectory" ;
        :references = "More information can be found at http://oceanobservatories.org/" ;
        :Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
        :date_created = "2016-06-14T16:07:44.374164" ;
        :id = "CP05MOAS-GL340-03-CTDGVM000-telemetered-ctdgv_m_glider_instrument" ;
        :requestUUID = "80a2377a-033b-4a1e-800d-2b3cfcd181cd" ;
        :contributor_role = "" ;
        :summary = "Dataset Generated by Stream Engine from Ocean Observatories Initiative" ;
        :keywords_vocabulary = "" ;
        :institution = "Ocean Observatories Initiative" ;
        :naming_authority = "org.oceanobservatories" ;
        :feature_Type = "point" ;
        :infoUrl = "http://oceanobservatories.org/" ;
        :license = "" ;
        :contributor_name = "" ;
        :uuid = "80a2377a-033b-4a1e-800d-2b3cfcd181cd" ;
        :creator_name = "Ocean Observatories Initiative" ;
        :title = "Data produced by Stream Engine version 1.0.1 for CP05MOAS-GL340-03-CTDGVM000-telemetered-ctdgv_m_glider_instrument" ;
        :sensor = "03-CTDGVM000" ;
        :standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention Standard Name Table 29" ;
        :acknowledgement = "" ;
        :project = "Ocean Observatories Initiative" ;
        :source = "CP05MOAS-GL340-03-CTDGVM000-telemetered-ctdgv_m_glider_instrument" ;
        :publisher_url = "http://oceanobservatories.org/" ;
        :creator_url = "http://oceanobservatories.org/" ;
        :nodc_template_version = "NODC_NetCDF_TimeSeries_Orthogonal_Template_v1.1" ;
        :subsite = "CP05MOAS" ;
        :processing_level = "L2" ;
        :time_coverage_resolution = "P69.19S" ;
        :geospatial_vertical_units = "meters" ;
        :geospatial_vertical_resolution = 0.1 ;
        :geospatial_vertical_positive = "down" ;
        :time_coverage_start = "2014-06-03T21:07:00.901Z" ;
        :time_coverage_end = "2014-06-03T22:58:45.412Z" ;
        :geospatial_lat_min = 40.049877166748 ;
        :geospatial_lat_max = 40.0509534606934 ;
        :geospatial_lon_min = -70.7527084350586 ;
        :geospatial_lon_max = -70.7489618530273 ;
        :DODS.strlen = 36 ;
        :DODS.dimName = "string36" ;
        :DODS_EXTRA.Unlimited_Dimension = "obs" ;
}
