netcdf illegal-vertical {
dimensions:
    time = 2;
variables:
    double time(time);
        time:standard_name = "time";
        time:units = "seconds since 1970-01-01";
    double z;
        z:long_name = "vertical position";
        z:axis = "Z";
        // units are missing
    double temp(time);
        temp:standard_name = "air_temperature";
        temp:units = "deg_C";

}
