netcdf sss_rc201401.v3.0cap {
dimensions:
	idlon = 360 ;
	idlat = 180 ;
variables:
	float idlon(idlon) ;
		idlon:long_name = "longitude" ;
		idlon:standard_name = "longitude" ;
		idlon:units = "degrees_east" ;
		idlon:comment = "midpoint of interval on uniform grid from -180 to 180 in 1 degree longitude increments" ;
		idlon:point_spacing = "1deg" ;
		idlon:axis = "X" ;
	float idlat(idlat) ;
		idlat:long_name = "latitude" ;
		idlat:standard_name = "latitude" ;
		idlat:units = "degrees_north" ;
		idlat:comment = "midpoint of interval on uniform grid from -90 to 90 in 1 degree latitude increments" ;
		idlat:point_spacing = "1deg" ;
		idlat:axis = "Y" ;
	float sss_cap(idlat, idlon) ;
		sss_cap:long_name = "Sea Surface Salinity" ;
		sss_cap:standard_name = "sea_surface_salinity" ;
		sss_cap:units = "1e-3" ;
		sss_cap:valid_min = 0.f ;
		sss_cap:valid_max = 45.f ;
		sss_cap:scale_factor = 1.f ;
		sss_cap:add_offset = 0.f ;
		sss_cap:grid_mapping = "Equirectangular" ;
		sss_cap:comment = "level-3 analysed sea surface salinity values obtained from the Combined Active Passive -CAP- algorithm with Rain Correction. Cell values are means for the temporal interval & 1degree spatial grid" ;
		sss_cap:_FillValue = -9999.f ;
		sss_cap:coordinates = "idlat idlon" ;
	char Equirectangular ;
		Equirectangular:grid_mapping_name = "latitude_longitude" ;
		Equirectangular:Standard_Parallel = 0.f ;
		Equirectangular:Longitude_of_Central_Meridian = 0.f ;
		Equirectangular:false_northing = 0.f ;
		Equirectangular:false_easting = 0.f ;
		Equirectangular:comment = "projection also referred to as Equidistant Cylindrical" ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:title = "Aquarius CAP 1x1 Deg Gridded Averaged Maps" ;
		:history = "DATA_SOURCE_VERSION 3.0" ;
		:institution = "JPL" ;
		:processing_level = "3" ;
		:cdm_data_type = "Grid" ;
		:date_issued = "2014-06-27T01:04:22Z" ;
		:date_created = "2014-06-27T01:04:22Z" ;
		:time_coverage_start = "01-2014" ;
		:time_coverage_end = "01-2014" ;
		:geospatial_lat_max = 90.f ;
		:geospatial_lat_min = -90.f ;
		:geospatial_lon_max = 180.f ;
		:geospatial_lon_min = -180.f ;
		:geospatial_lat_resolution = 1.f ;
		:geospatial_lon_resolution = 1.f ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:platform = "Aquarius/SAC-D" ;
		:sensor = "Aquarius" ;
		:project = "Aquarius" ;
		:product_version = "3.0" ;
		:keywords_vocabulary = "http://gcmd.gsfc.nasa.gov/Resources/valids/gcmd_parameters.html" ;
		:keywords = "SURFACE SALINITY, SALINITY, AQUARIUS, Jet Propulsion Laboratory, NASA, http://aquarius.nasa.gov/, AQUARIUS SAC-D, Aquarius Scatterometer, Aquarius Radiometer" ;
		:summary = "Version 3.0 Aquarius CAP Level 3 products contain mapped Aquarius sea surface salinity or wind speed data based on the Combined Active Passive (CAP) algorithm. CAP is a P.I. produced data set developed and provided by the JPL Climate Oceans and Solid Earth section.  (For further details see   http://podaac.jpl.nasa.gov/dataset/AQUARIUS_L3_SSS_CAP_7DAY_V3 )" ;
		:creator_name = "Simon H. Yueh" ;
		:creator_email = "Simon.H.Yueh@jpl.nasa.gov" ;
		:creator_url = "http://science.jpl.nasa.gov/COSE/index.cfm" ;
		:publisher_name = "Simon H. Yueh" ;
		:publisher_email = "Simon.H.Yueh@jpl.nasa.gov" ;
		:publisher_url = "http://science.jpl.nasa.gov/COSE/index.cfm" ;
		:contributor_name = "Wenqing Tang, Alex Fore, Akiko Hayashi" ;
		:contributor_role = "Aquarius-CAP algorithm geophysical model functions, CAP algorithm operational setup and L2 processing, L3 algorithm implementation, processing and data staging " ;
		:Data_Type = "1x1 Deg Gridded Bin Averaged Maps" ;
		:VARIABLE_1 = "sss_cap(nlon,nlat)" ;
		:First_Index = "Longitude" ;
		:Second_Index = "Latitude" ;
		:Map_Time_Range = "201401" ;
		:Search_Radius_KM = "      111.000" ;
		:Half_Power_Point_KM = "      75.0000" ;
		:Binning_Method = "Gaussian" ;
		:Land_Fraction = "    0.0100000" ;
		:Ice_Fraction = "  0.000500000" ;
		:Minimum_Bin_Pts = "      10.0000" ;
		:VARIABLE_2 = "ice_frac(nlon,nlat)" ;
}
