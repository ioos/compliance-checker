netcdf rhgrid {
dimensions:
	londim = 128 ;
	latdim = 64 ;
	rgrid = 6144 ;
variables:
	float PS(rgrid) ;
		PS:long_name = "surface pressure" ;
		PS:units = "Pa" ;
		PS:coordinates = "lon lat" ;
	float lon(rgrid) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
	float lat(rgrid) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
	float rgrid(rgrid) ;
		rgrid:compress = "latdim londim" ;
}
