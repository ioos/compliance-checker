netcdf conv_multi {

// global attributes:
		:featureType = "timeSeries" ;
		:NCO = "4.4.2" ;
		:history = "Wed Feb 25 15:10:07 2015: ncatted -a Conventions,global,o,c,CF-1.6 ,ACDD awfu.nc\nWed Feb 25 15:09:40 2015: ncks -x -v lat,lon,time,height,water_temp compliance_checker/tests/data/example-grid.nc awfu.nc" ;
		:Conventions = "CF-1.6 ,ACDD" ;
}
