netcdf forecast_reference.cdl {
dimensions:
    time = 2 ;
    lat = 4 ;
    lon = 4 ;
variables:
    float time(time) ;
        time:units = "seconds since 1970-01-01" ;
        time:standard_name = "time" ;
        time:calendar = "gregorian" ;
        time:axis = "T" ;
    float lat(lat) ;
        lat:units = "degrees_north" ;
        lat:standard_name = "latitude" ;
        lat:axis = "Y" ;
    float lon(lon) ;
        lon:units = "degrees_east" ;
        lon:standard_name = "longitude" ;
        lon:axis = "X" ;
    float air_temp(time, lon, lat) ;
        air_temp:units = "deg_C" ;
        air_temp:standard_name = "air_temperature";
    float forecast_reference_time(time) ;
        forecast_reference_time:units = "seconds since 1970-01-01" ;
        forecast_reference_time:standard_name = "forecast_reference_time" ;
    float forecast_hour(time) ;
        forecast_hour:units = "hours" ;
        forecast_hour:standard_name = "forecast_period" ;

    :featureType = "grid" ;

}
