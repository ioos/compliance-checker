netcdf timeseries-orthogonal {
dimensions:
 station = 10 ;  // measurement locations
 name_strlen = 12;
 time = UNLIMITED ;
variables:
    float humidity(time, station) ;
        humidity:standard_name = "specific_humidity" ;
        humidity:coordinates = "lat lon alt" ;
    double time(time) ;
        time:standard_name = "time";
        time:long_name = "time of measurement" ;
        time:units = "days since 1970-01-01 00:00:00" ;
    float lon(station) ;
        lon:standard_name = "longitude";
        lon:long_name = "station longitude";
        lon:units = "degrees_east";
    float lat(station) ;
        lat:standard_name = "latitude";
        lat:long_name = "station latitude" ;
        lat:units = "degrees_north" ;
    float alt(station) ;
        alt:long_name = "vertical distance above the surface" ;
        alt:standard_name = "height" ;
        alt:units = "m";
        alt:positive = "up";
        alt:axis = "Z";
    char station_name(station, name_strlen) ;
        station_name:long_name = "station name" ;
        station_name:cf_role = "timeseries_id";
// attributes
    :featureType = "timeSeries";
    :Conventions = "CF-1.6";
    :institution = "CF";
    :source = "fake";
    :references = "http://cfconventions.org/cf-conventions/v1.6.0/cf-conventions.html#_point_data";
    :title = "CF-1.6 H.2.1 Orthogonal multidimensional array representation of time series";
    :history = "2016-10-31T18:32Z - File Created";

}
