netcdf time_units {
dimensions:
    time = 10 ;
variables:
    uint64 time(time) ;
        time:units = "seconds since 1970-01-01" ;
        time:standard_name = "time" ;
        time:calendar = "gregorian" ;
    float temperature(time) ;
        temperature:units = "days since 1970-01-01" ;
        temperature:standard_name = "sea_water_temperature" ;

// global attributes:
		:featureType = "timeSeries" ;
}

