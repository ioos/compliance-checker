netcdf vertical_coords {
dimensions:
    time = 2;
variables:
    double time(time);
        time:units = "seconds since 1970-01-01";
        time:standard_name = "time";
        time:axis = "T";
    // height is not a coordinate variable, does not define a standard name, or
    // axis but is referenced by coordinates, this is a valid cf auxiliary
    // coordinate.
    float height(time);
        height:units = "hPa";
    float temperature(time);
        temperature:standard_name = "air_temperature";
        temperature:units = "deg_C";
        temperature:coordinates = "time height lat lon";
    :title = "Example dataset defining vertical coordinates";
    :institution = "IOOS";
    :source = "imagination";
    :history = "2016-10-24T17:00Z - Created";
    :references = "CF 1.6";

}
