netcdf rotated_pole_grid {
dimensions:
    rlon = 2;
    rlat = 2;
    lev = 2;
variables:
    float temperature(lev, rlat, rlon);
        temperature:long_name = "temperature";
        temperature:standard_name = "air_temperature";
        temperature:units = "K";
        temperature:coordinates = "lon lat";
        temperature:grid_mapping = "rotated_pole";

    char rotated_pole;
        rotated_pole:grid_mapping_name = "rotated_latitude_longitude";
        rotated_pole:grid_north_pole_latitude = 32.5;
        rotated_pole:grid_north_pole_longitude = 170.;
    float rlon(rlon);
        rlon:long_name = "longitude in rotated pole grid";
        rlon:units = "degrees";
        rlon:standard_name = "grid_longitude";
        rlon:axis = "X";

    float rlat(rlat);
        rlat:long_name = "latitude in rotated pole grid";
        rlat:units = "degrees";
        rlat:standard_name = "grid_latitude";
        rlat:axis = "Y";

    float lev(lev);
        lev:long_name = "pressure level";
        lev:units = "hPa";
        lev:axis = "Z";

    float lon(rlat, rlon);
        lon:long_name = "longitude";
        lon:units = "degrees_east";
        lon:standard_name = "longitude";

    float lat(rlat, rlon);
        lat:long_name = "latitude";
        lat:units = "degrees_north";
        lat:standard_name = "latitude";

}
