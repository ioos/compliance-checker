netcdf bad_data_type {
dimensions:
	time = 3 ;
	latitude = 1 ;
	longitude = 1 ;
	power = 1 ;
variables:
	double time(time) ;
	double latitude(latitude) ;
		latitude:units = "Degrees_N" ;
		latitude:axis = "Y" ;
		latitude:bounds = "salinity" ;
	double longitude(longitude) ;
		longitude:units = "Degrees_E" ;
		longitude:compress = "longitude latitude" ;
	int64 temp(time, time) ;
		temp:_FillValue = -999L ;
		temp:valid_min = 0L ;
		temp:valid_max = 10L ;
		temp:units = "K" ;
		temp:add_offset = "c" ;
		temp:scale_factor = 5L ;
		temp:compress = "time longitudeZZ" ;
	double salinity(latitude, longitude, time) ;
		salinity:_FillValue = 1. ;
		salinity:valid_min = -10L ;
		salinity:valid_max = 10L ;
		salinity:institution = 10L ;
		salinity:units = "Chad Pennington" ;
		salinity:standard_name = "Chadwick Penington" ;
		salinity:axis = "Time" ;
		salinity:coordinates = "latitude longitudeZZ time" ;
		salinity:add_offset = 5. ;
		salinity:scale_factor = 5. ;
	double longitudeZZ(longitude) ;
		longitudeZZ:_FillValue = 1. ;
		longitudeZZ:coordinates = "longitude" ;
	double really_bad(latitude, power) ;

// global attributes:
		:featureType = "pointzz" ;
data:

 time = _, _, _ ;

 latitude = _ ;

 longitude = _ ;

 temp =
  _, _, _,
  _, _, _,
  _, _, _ ;

 salinity =
  _, _, _ ;

 longitudeZZ = _ ;

 really_bad =
  _ ;
}

