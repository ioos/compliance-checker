netcdf bad_region {
dimensions:
	time = 3 ; // (3 currently)
	strlen = 14 ;
	latitude = 1 ;
	longitude = 1 ;
variables:
	double time(time) ;
	double latitude(latitude) ;
		latitude:units = "Degrees_N" ;
		latitude:axis = "Y" ;
	double longitude(longitude) ;
		longitude:units = "Degrees_E" ;
    double temp(time);
		temp:units = "K" ;
	double salinity(latitude, longitude, time) ;
		salinity:_FillValue = 1. ;
		salinity:valid_min = -10L ;
		salinity:valid_max = 10L ;
		salinity:institution = 10L ;
		salinity:units = "Chad Pennington" ;
		salinity:standard_name = "Chadwick Penington" ;
		salinity:axis = "Time" ;
		salinity:coordinates = "latitude longitudeZZ time" ;
	double longitudeZZ(longitude) ;
		longitudeZZ:_FillValue = 1. ;
	char neverland(strlen) ;
		neverland:standard_name = "region" ;
	char geo_region(strlen) ;
		geo_region:standard_name = "region" ;
data:

 time = 1., 2., 3. ;

 latitude = 40. ;

 longitude = -60. ;

 temp = _, _, _;

 salinity = 0.65873145682807, 0.715646913770724, _ ;

 longitudeZZ = _ ;

 neverland = "Neverland" ;

 geo_region = "Atlantic_Ocean" ;
}
