netcdf ints64 {
dimensions:
    time = 10 ;
variables:
    uint64 time(time) ;
        time:units = "seconds since 1970-01-01" ;
        time:standard_name = "time" ;
        time:calendar = "gregorian" ;
    uint64 temp_counts(time) ;
        temp_counts:units = "1" ;

// global attributes:
		:featureType = "timeSeries" ;
data:

time = 1406689200, 1406692800, 1406696400, 1406700000, 1406703600 ;
temp_counts = 1, 2, 3, 4, 5 ;
}
