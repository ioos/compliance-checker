netcdf timeseries-profile-single-station {
dimensions:
    time = 2;
    z = 10;
variables:
    double time(time);
        time:standard_name = "time";
        time:long_name = "Time";
        time:axis = "T";
        time:units = "seconds since 1970-01-01T00:00:00Z";
    float lat;
        lat:standard_name = "latitude";
        lat:units = "degrees_north";
        lat:axis = "Y";
        lat:long_name = "Latitude";
    float lon;
        lon:standard_name = "longitude";
        lon:units = "degrees_east";
        lon:axis = "X";
        lon:long_name = "Longitude";
    float z(z);
        z:standard_name = "depth";
        z:positive = "down";
        z:units = "m";
        z:long_name = "Depth below surface";

    float temperature(time, z);
        temperature:standard_name = "sea_water_temperature";
        temperature:units = "deg_C";
        temperature:long_name = "Seawater Temperature";
        temperature:coordinates = "time lat lon z";

}




