netcdf \2dim-grid {
dimensions:
	lev = 5 ;
	yc = 2 ;
	xc = 2 ;
variables:
	float T(lev, yc, xc) ;
		T:long_name = "temperature" ;
		T:units = "K" ;
		T:coordinates = "lon lat" ;
	float xc(xc) ;
		xc:axis = "X" ;
		xc:long_name = "x-coordinate in Cartesian system" ;
		xc:units = "m" ;
	float yc(yc) ;
		yc:axis = "Y" ;
		yc:long_name = "y-coordinate in Cartesian system" ;
		yc:units = "m" ;
	float lev(lev) ;
		lev:long_name = "pressure level" ;
		lev:units = "hPa" ;
	float lon(yc, xc) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
	float lat(yc, xc) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
	float quality_control(yc, xc) ;
		quality_control:long_name = "quality control" ;
		quality_control:flag_meanings = "flag meanings" ;
data:

 T =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _ ;

 xc = _, _ ;

 yc = _, _ ;

 lev = _, _, _, _, _ ;

 lon =
  _, _,
  _, _ ;

 lat =
  _, _,
  _, _ ;

 quality_control =
  _, _,
  _, _ ;
}
