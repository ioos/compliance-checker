netcdf sea_water_temperature {
dimensions:
    maxStrlen64 = 64 ;
    time = 14 ;
variables:
    char feature_type_instance(maxStrlen64) ;
        feature_type_instance:cf_role = "timeseries_id" ;
        feature_type_instance:long_name = "Identifier for each feature type instance" ;
    double latitude ;
        latitude:units = "degrees_north" ;
        latitude:standard_name = "latitude" ;
        latitude:long_name = "sensor latitude" ;
    double longitude ;
        longitude:units = "degrees_east" ;
        longitude:standard_name = "longitude" ;
        longitude:long_name = "sensor longitude" ;
    int crs ;
        crs:long_name = "http://www.opengis.net/def/crs/EPSG/0/4326" ;
        crs:grid_mapping_name = "latitude_longitude" ;
        crs:epsg_code = "EPSG:4326" ;
        crs:semi_major_axis = 6378137. ;
        crs:inverse_flattening = 298.257223563 ;
    int platform ;
        platform:definition = "http://mmisw.org/ont/ioos/definition/stationID" ;
        platform:short_name = "kibesillah_hill_intertidal_shore_station" ;
        platform:long_name = "urn:ioos:station:cencoos:kibesillah_hill_intertidal_shore_station" ;
        platform:ioos_code = "urn:ioos:station:cencoos:kibesillah_hill_intertidal_shore_station" ;
    int time(time) ;
        time:units = "seconds since 1970-01-01T00:00:00Z" ;
        time:standard_name = "time" ;
        time:long_name = "time of measurement" ;
        time:calendar = "gregorian" ;
    double height ;
        height:_FillValue = -9999.9 ;
        height:grid_mapping = "crs" ;
        height:long_name = "height of the sensor relative to the water surface" ;
        height:standard_name = "depth" ;
        height:positive = "down" ;
        height:units = "m" ;
        height:axis = "Z" ;
    double sea_water_temperature(time) ;
        sea_water_temperature:instrument = "sea_water_temperature_instrument" ;
        sea_water_temperature:coordinates = "time height latitude longitude" ;
        sea_water_temperature:standard_name = "sea_water_temperature" ;
        sea_water_temperature:units = "degree_Celsius" ;
        sea_water_temperature:grid_mapping = "crs" ;
        sea_water_temperature:platform = "platform" ;
        sea_water_temperature:_FillValue = -9999.9 ;
    int sea_water_temperature_instrument ;
        sea_water_temperature_instrument:ioos_code = "urn:ioos:sensor:cencoos:kibesillah_hill_intertidal_shore_station:sea_water_temperature" ;
        sea_water_temperature_instrument:short_name = "sea_water_temperature" ;
        sea_water_temperature_instrument:definition = "http://mmisw.org/ont/ioos/definition/sensorID" ;
        sea_water_temperature_instrument:long_name = "urn:ioos:sensor:cencoos:kibesillah_hill_intertidal_shore_station:sea_water_temperature" ;

// global attributes:
        :contributor_role = "Data Provider" ;
        :creator_url = "http://cencoos.org/" ;
        :creator_type = "institution" ;
        :contributor_name = "Central & Northern California Ocean Observing System (CeNCOOS)" ;
        :commment = "This is an aggregation of the entire archive available for this platform and variable and is updated every three days for live data streams. It may not include quasi real-time data." ;
        :license = "The data may be used and redistributed for free but is not intended for legal use, since it may contain inaccuracies. No person or group associated with this data makes any warranty, express or implied, including warranties of merchantability and fitness for a particular purpose, or assumes any legal liability for the accuracy, completeness, or usefulness, of this information." ;
        :publisher_email = "axiom+archives@axiomdatascience.com" ;
        :institution = "Central & Northern California Ocean Observing System (CeNCOOS)" ;
        :creator_email = "jpatterson@mbari.org" ;
        :keywords_vocabulary = "GCMD Science Keywords" ;
        :creator_name = "Central & Northern California Ocean Observing System (CeNCOOS)" ;
        :processing_level = "Raw data stream, no quality checks performed" ;
        :publisher_name = "Axiom Data Science" ;
        :naming_authority = "cencoos" ;
        :description = "Full set of archive data from Kibesillah Hill Intertidal Shore Station" ;
        :publisher_url = "http://axiomdatascience.com" ;
        :summary = "Kibesillah Hill Intertidal Shore Station" ;
        :keywords = "In Situ Ocean-based platforms, Oceans" ;
        :id = "kibesillah_hill_intertidal_shore_station" ;
        :standard_name_vocabulary = "CF Standard Name Table v25" ;
        :Conventions = "CF-1.6" ;
        :Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
        :date_created = "2016-07-16T22:46:00Z" ;
        :date_issued = "2016-07-16T22:46:00Z" ;
        :cdm_data_type = "Station" ;
        :history = "Created by Axiom NetCDF Archiver\n",
            "2016-07-16T22:46:00Z - pyaxiom - File created using pyaxiom" ;
        :geospatial_lat_min = 39.6004 ;
        :geospatial_lat_max = 39.6004 ;
        :geospatial_lat_units = "degrees_north" ;
        :geospatial_lon_min = -123.7892 ;
        :geospatial_lon_max = -123.7892 ;
        :geospatial_lon_units = "degrees_east" ;
        :platform = "platform" ;
        :time_coverage_start = "2009-01-01T08:00:00" ;
        :time_coverage_end = "2015-12-29T13:19:59" ;
        :time_coverage_duration = "P220598399S" ;
        :time_coverage_resolution = "P599S" ;
        :geospatial_vertical_units = "meters" ;
        :geospatial_vertical_positive = "down" ;
        :featureType = "timeSeries" ;
        :geospatial_vertical_resolution = "0" ;
        :geospatial_vertical_min = 0.1524 ;
        :geospatial_vertical_max = 0.1524 ;
        :DODS.strlen = 65 ;
        :DODS.dimName = "feature_type_instance" ;
}
