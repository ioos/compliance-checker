netcdf Hurricane_Ike_2D_preliminary_run_1_without_waves {
dimensions:
    Layer = 1 ;
    LayerInterf = 2 ;
    bounds4 = 4 ;
    grid_m = 4 ;
    grid_n = 4 ;
    m = 4 ;
    n = 4 ;
    time = 8 ;
    time_bounds = 2 ;
variables:
    double time(time) ;
        time:standard_name = "time" ;
        time:long_name = "time" ;
        time:units = "days since 1970-01-01 00:00:00 " ;
        time:axis = "T" ;
        time:delft3d_name = "map-info-series:ITMAPC map-const:ITDATE map-const:DT map-const:TUNIT" ;
        time:actual_range = 14131., 14136.25 ;
    double time_bounds(time_bounds, time) ;
        time_bounds:long_name = "time bounds" ;
        time_bounds:actual_range = "2008-09-09 00:00:00\t2008-09-14 06:00:00" ;
    float longitude(m, n) ;
        longitude:standard_name = "longitude" ;
        longitude:long_name = "grid cell centers, longitude-coordinate" ;
        longitude:units = "degrees_east" ;
        longitude:axis = "X" ;
        longitude:_FillValue = NaNf ;
        longitude:missing_value = NaNf ;
        longitude:actual_range = -97.8499984741211, -80.25 ;
        longitude:delft3d_name = "map-const:XZ map-const:KCS map-const:CODW map-const:COORDINATES" ;
    float latitude(m, n) ;
        latitude:standard_name = "latitude" ;
        latitude:long_name = "grid cell centers, latitude-coordinate" ;
        latitude:units = "degrees_north" ;
        latitude:axis = "Y" ;
        latitude:_FillValue = NaNf ;
        latitude:missing_value = NaNf ;
        latitude:actual_range = 18.1499996185303, 30.75 ;
        latitude:delft3d_name = "map-const:YZ map-const:KCS map-const:YWAT map-const:CODW map-const:COORDINATES" ;
    float grid_longitude(m, n, bounds4) ;
        grid_longitude:long_name = "grid cell corners, longitude-bounds" ;
        grid_longitude:units = "degrees_east" ;
        grid_longitude:_FillValue = NaNf ;
        grid_longitude:missing_value = NaNf ;
        grid_longitude:actual_range = -97.9000015258789, 0. ;
        grid_longitude:delft3d_name = "map-const:XCOR map-const:CODB map-const:COORDINATES" ;
    float grid_latitude(m, n, bounds4) ;
        grid_latitude:long_name = "grid cell corners, latitude-bounds" ;
        grid_latitude:units = "degrees_north" ;
        grid_latitude:_FillValue = NaNf ;
        grid_latitude:missing_value = NaNf ;
        grid_latitude:actual_range = 0., 30.7999992370605 ;
        grid_latitude:delft3d_name = "map-const:YCOR map-const:CODB map-const:COORDINATES" ;
    float k(Layer) ;
        k:long_name = "layer index" ;
        k:units = "1" ;
        k:axis = "Z" ;
        k:comment = "The surface layer has index k=1, the bottom layer has index kmax." ;
        k:delft3d_name = "map-const:KMAX map-const:LAYER_MODEL" ;
    float Layer(Layer) ;
        Layer:long_name = "sigma at layer midpoints" ;
        Layer:standard_name = "ocean_sigma_coordinate" ;
        Layer:positive = "up" ;
        Layer:formula_terms = "sigma: Layer eta: waterlevel depth: depth" ;
        Layer:actual_range = -0.5, -0.5 ;
        Layer:comment = "The surface layer has index k=1 and is sigma=0, the bottom layer has index kmax and is sigma=-1." ;
        Layer:delft3d_name = "map-const:KMAX map-const:LAYER_MODEL map-const:THICK" ;
    float LayerInterf(LayerInterf) ;
        LayerInterf:long_name = "sigma at layer interfaces" ;
        LayerInterf:standard_name = "ocean_sigma_coordinate" ;
        LayerInterf:positive = "up" ;
        LayerInterf:formula_terms = "sigma: LayerInterf eta: waterlevel depth: depth" ;
        LayerInterf:actual_range = -1., 0. ;
        LayerInterf:comment = "The surface layer has index k=1 and is sigma=0, the bottom layer has index kmax and is sigma=-1." ;
        LayerInterf:delft3d_name = "map-const:KMAX map-const:LAYER_MODEL map-const:THICK" ;
    float grid_depth(grid_m, grid_n) ;
        grid_depth:standard_name = "sea_floor_depth_below_sea_level" ;
        grid_depth:long_name = "depth of cell corners" ;
        grid_depth:units = "m" ;
        grid_depth:_FillValue = NaNf ;
        grid_depth:missing_value = NaNf ;
        grid_depth:actual_range = NaN, NaN ;
        grid_depth:delft3d_name = "map-const:DP map-const:DP0 map-const:DPS map-const:DRYFLP" ;
        grid_depth:comment = "" ;
    float depth(m, n) ;
        depth:standard_name = "sea_floor_depth_below_sea_level" ;
        depth:long_name = "depth of cell centers" ;
        depth:units = "m" ;
        depth:coordinates = "latitude longitude" ;
        depth:_FillValue = NaNf ;
        depth:missing_value = NaNf ;
        depth:actual_range = -7146.62353515625, 67.0625 ;
        depth:delft3d_name = "map-const:DPS0 map-const:KCS" ;
        depth:comment = "" ;
    float zactive(m, n) ;
        zactive:long_name = "active water-level point" ;
        zactive:units = "1" ;
        zactive:coordinates = "latitude longitude" ;
        zactive:_FillValue = NaNf ;
        zactive:missing_value = NaNf ;
        zactive:actual_range = 0., 1. ;
        zactive:delft3d_name = "map-const:KCS" ;
    float area(m, n) ;
        area:standard_name = "cell_area" ;
        area:long_name = "area of grid cells" ;
        area:units = "degrees2" ;
        area:coordinates = "latitude longitude" ;
        area:_FillValue = NaNf ;
        area:missing_value = NaNf ;
        area:actual_range = 0.00999969482654706, 0.0100006485008635 ;
        area:delft3d_name = "map-const:GSQS map-const:KCS" ;
        area:comment = "This is the exact area spanned geometrically by the 4 corner points. This is not identical to the area GSQS used internally in Delft3D for mass-conservation!" ;
    float waterlevel(time, m, n) ;
        waterlevel:standard_name = "sea_surface_height_above_geoid" ;
        waterlevel:long_name = "water level" ;
        waterlevel:units = "m" ;
        waterlevel:coordinates = "latitude longitude" ;
        waterlevel:_FillValue = NaNf ;
        waterlevel:missing_value = NaNf ;
        waterlevel:actual_range = -2.13350892066956, 67.0625 ;
        waterlevel:cell_methods = "time: point             " ;
        waterlevel:delft3d_name = "map-series:S1 map-const:KCS" ;
    float velocity_x(time, Layer, m, n) ;
        velocity_x:standard_name = "eastward_sea_water_velocity" ;
        velocity_x:long_name = "velocity, lon-component" ;
        velocity_x:units = "m/s" ;
        velocity_x:coordinates = "latitude longitude" ;
        velocity_x:_FillValue = NaNf ;
        velocity_x:missing_value = NaNf ;
        velocity_x:actual_range = -2.64120197296143, 1.0327941775322 ;
        velocity_x:cell_methods = "time: point             " ;
        velocity_x:delft3d_name = "map-series:U1 map-series:V1 map-const:ALFAS map-const:KCU map-const:KCV map-const:KFU map-const:KFV map-const:KCS" ;
    float velocity_y(time, Layer, m, n) ;
        velocity_y:standard_name = "northward_sea_water_velocity" ;
        velocity_y:long_name = "velocity, lat-component" ;
        velocity_y:units = "m/s" ;
        velocity_y:coordinates = "latitude longitude" ;
        velocity_y:_FillValue = NaNf ;
        velocity_y:missing_value = NaNf ;
        velocity_y:actual_range = -1.52386540174484, 6.19752788543701 ;
        velocity_y:cell_methods = "time: point             " ;
        velocity_y:delft3d_name = "map-series:U1 map-series:V1 map-const:ALFAS map-const:KCU map-const:KCV map-const:KFU map-const:KFV map-const:KCS" ;
    float tau_x(time, m, n) ;
        tau_x:standard_name = "surface_downward_northward_stress" ;
        tau_x:long_name = "bed shear stress, x-component" ;
        tau_x:units = "N/m2" ;
        tau_x:coordinates = "latitude longitude" ;
        tau_x:_FillValue = NaNf ;
        tau_x:missing_value = NaNf ;
        tau_x:actual_range = -93.8008499145508, 157.384719848633 ;
        tau_x:cell_methods = "time: point             " ;
        tau_x:delft3d_name = "map-series:TAUKSI map-const:TAUETA map-const:ALFAS map-const:KCS" ;
    float tau_y(time, m, n) ;
        tau_y:standard_name = "surface_downward_eastward_stress" ;
        tau_y:long_name = "bed shear stress, y-component" ;
        tau_y:units = "N/m2" ;
        tau_y:coordinates = "latitude longitude" ;
        tau_y:_FillValue = NaNf ;
        tau_y:missing_value = NaNf ;
        tau_y:actual_range = -2561.92041015625, 373.899017333984 ;
        tau_y:cell_methods = "time: point             " ;
        tau_y:delft3d_name = "map-series:TAUKSI map-const:TAUETA map-const:ALFAS map-const:KCS" ;

// global attributes:
        :title = "Pr Inundation Tropical : NRL : DELFT3D : Hurricane Ike 2D preliminary run 1 without waves" ;
        :institution = "" ;
        :source = "Delft3D trim file" ;
        :history = "Original filename: trim-ike.dat, Deltares, FLOW2D3D Version 5.01.00.2350, Mar 13 2013, 15:39:06, file version: 3.54.29, file date:2013-04-04 15:21:00, transformation to netCDF: $HeadURL: https://svn.oss.deltares.nl/repos/openearthtools/trunk/matlab/applications/delft3d/vs_trim2nc.m $ $Id: vs_trim2nc.m 10615 2014-04-28 10:03:00Z boer_g $" ;
        :references = "http://svn.oss.deltares.nl" ;
        :email = "" ;
        :comment = "" ;
        :version = "Deltares, FLOW2D3D Version 5.01.00.2350, Mar 13 2013, 15:39:06, file version: 3.54.29" ;
        :Conventions = "CF-1.6" ;
        :terms_for_use = "These data can be used freely for research purposes provided that the following source is acknowledged: " ;
        :disclaimer = "This data is made available in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE." ;
        :delft3d_description = "                              \n",
            "                              \n",
            "                              \n",
            "                              \n",
            "                              \n",
            "                              \n",
            "                              \n",
            "                              \n",
            "                              \n",
            "                              \n",
            "" ;
        :time_coverage_start = "2008-09-09T00:00" ;
        :time_coverage_end = "2008-09-14T06:00" ;
        :geospatial_lat_min = 18.1499996185303 ;
        :geospatial_lat_max = 30.75 ;
        :geospatial_lat_units = "dergees_north" ;
        :geospatial_lon_min = -97.8499984741211 ;
        :geospatial_lon_max = -80.25 ;
        :geospatial_lon_units = "dergees_east" ;
        :geospatial_vertical_min = -67.0625 ;
        :geospatial_vertical_max = 7146.62353515625 ;
        :geospatial_vertical_units = "m" ;
        :geospatial_vertical_positive = "down" ;
        :id = "pr_inundation_tropical.NRL_DELFT3D.Hurricane_Ike_2D_preliminary_run_1_without_waves" ;
        :cdm_data_type = "" ;
        :summary = "A test of Hurricane Ike (2008) using Delft3D" ;
        :ncmlFile = "/data/comt_2/pr_inundation_tropical/NRL_Delft3D/Hurricane_Ike_2D_preliminary_run_1_without_waves/00_dir.ncml" ;
}
