netcdf string_type_variable {
dimensions:
        lon = 10 ;
variables:
        double lon(lon) ;
		lon:long_name = "location of something a specific longitudinal coordinates" ;
		lon:axis = "X" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
        string j(lon) ;
		j:long_name = "name of each measurement location" ;

// global attributes:
	:Conventions = "CF-1.7" ;
	:title = "file to test proper processing of string-type variables" ;
	:history = "2020-07-22T17:04: hand-made" ;
}

