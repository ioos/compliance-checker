
netcdf SWAN_Tutuila_Regional_Wave_Model_best {
dimensions:
	lat = 4 ;
	lon = 4 ;
	time = 8 ;
	z = 1 ;
variables:
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:short_name = "lon" ;
		lon:axis = "x" ;
		lon:_CoordinateAxisType = "Lon" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:short_name = "lat" ;
		lat:axis = "y" ;
		lat:_CoordinateAxisType = "Lat" ;
	float z(z) ;
		z:units = "meters" ;
		z:long_name = "depth below mean sea level" ;
		z:standard_name = "depth" ;
		z:short_name = "depth" ;
		z:axis = "z" ;
		z:_CoordinateAxisType = "Height" ;
	double time(time) ;
		time:long_name = "Forecast time for ForecastModelRunCollection" ;
		time:standard_name = "time" ;
		time:calendar = "proleptic_gregorian" ;
		time:units = "hours since 2013-02-18 00:00:00.000 UTC" ;
		time:missing_value = NaN ;
		time:_CoordinateAxisType = "Time" ;
	double time_run(time) ;
		time_run:long_name = "run times for coordinate = time" ;
		time_run:standard_name = "forecast_reference_time" ;
		time_run:calendar = "proleptic_gregorian" ;
		time_run:units = "hours since 2013-02-18 00:00:00.000 UTC" ;
		time_run:missing_value = NaN ;
		time_run:_CoordinateAxisType = "RunTime" ;
	double time_offset(time) ;
		time_offset:long_name = "offset hour from start of run for coordinate = time" ;
		time_offset:standard_name = "forecast_period" ;
		time_offset:calendar = "proleptic_gregorian" ;
		time_offset:units = "hours since 2013-02-18T00:00:00Z" ;
		time_offset:missing_value = NaN ;
	float shgt(time, z, lat, lon) ;
		shgt:units = "meters" ;
		shgt:long_name = "significant wave height" ;
		shgt:standard_name = "sea_surface_wave_significant_height" ;
		shgt:short_name = "hs" ;
		shgt:valid_range = 0.f, 20.f ;
		shgt:_FillValue = NaNf ;
		shgt:coordinates = "time_run time z lat lon " ;
	float mper(time, z, lat, lon) ;
		mper:units = "seconds" ;
		mper:long_name = "mean wave period" ;
		mper:standard_name = "sea_surface_wave_mean_period_from_variance_spectral_density_second_frequency_moment" ;
		mper:short_name = "mper" ;
		mper:valid_range = 0.f, 30.f ;
		mper:_FillValue = NaNf ;
		mper:coordinates = "time_run time z lat lon " ;
	float mdir(time, z, lat, lon) ;
		mdir:units = "degrees" ;
		mdir:long_name = "mean wave direction" ;
		mdir:standard_name = "sea_surface_wave_from_direction" ;
		mdir:short_name = "mdir" ;
		mdir:valid_range = 0.f, 360.f ;
		mdir:_FillValue = NaNf ;
		mdir:coordinates = "time_run time z lat lon " ;
	float pper(time, z, lat, lon) ;
		pper:units = "seconds" ;
		pper:long_name = "peak wave period" ;
		pper:standard_name = "sea_surface_wave_period_at_variance_spectral_density_maximum" ;
		pper:short_name = "pper" ;
		pper:valid_range = 0.f, 30.f ;
		pper:_FillValue = NaNf ;
		pper:coordinates = "time_run time z lat lon " ;
	float pdir(time, z, lat, lon) ;
		pdir:units = "degrees" ;
		pdir:long_name = "peak wave direction" ;
		pdir:standard_name = "sea_surface_wave_from_direction" ;
		pdir:short_name = "pdir" ;
		pdir:valid_range = 0.f, 360.f ;
		pdir:_FillValue = NaNf ;
		pdir:coordinates = "time_run time z lat lon " ;

// global attributes:
		:title = "Simulating WAves Nearshore (SWAN) Regional Wave Model: Tutuila, American Samoa" ;
		:_CoordSysBuilder = "ucar.nc2.dataset.conv.CF1Convention" ;
		:Conventions = "Unidata Dataset Discovery v1.0, CF-1.4" ;
		:cdm_data_type = "Grid" ;
		:featureType = "GRID" ;
		:location = "Proto fmrc:SWAN_Tutuila_Regional_Wave_Model" ;
		:id = "swan_tutuila" ;
		:naming_authority = "org.pacioos" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0, CF-1.4" ;
		:Metadata_Link = "http://pacioos.org/metadata/swan_tutuila.html" ;
		:ISO_Topic_Categories = "oceans" ;
		:summary = "Simulating WAves Nearshore (SWAN) regional wave model 7-day output with a 5-day hourly forecast for the island of Tutuila, American Samoa at approximately 500-m resolution. This high-resolution model is utilized to capture shallow water effects and nearshore coastal dynamics such as refracting, shoaling, and smaller scale shadowing. It is run directly after the Samoa regional WaveWatch III (WW3) wave model has completed. Please note that this nested model setup is in the testing and validation phase. While considerable effort has been made to implement all model components in a thorough, correct, and accurate manner, numerous sources of error are possible. As such, please use these data with the caution appropriate for any ocean related activity." ;
		:keywords = "Earth Science Services > Models > Ocean General Circulation Models (OGCM)/Regional Ocean Models, Earth Science Services > Models > Weather Research/Forecast Models, Earth Science > Oceans > Ocean Waves > Significant Wave Height, Earth Science > Oceans > Ocean Waves > Wave Period, Earth Science > Oceans > Ocean Waves > Wave Speed/Direction" ;
		:keywords_vocabulary = "GCMD Science Keywords" ;
		:standard_name_vocabulary = "CF-1.4" ;
		:comment = "Model runs produced by Dr. Kwok Fai Cheung (cheung@hawaii.edu)." ;
		:geospatial_lat_min = -14.4 ;
		:geospatial_lat_max = -14.15 ;
		:geospatial_lon_min = 189. ;
		:geospatial_lon_max = 189.6 ;
		:geospatial_vertical_min = 0. ;
		:geospatial_vertical_max = 0. ;
		:time_coverage_start = "2013-02-18T21:00:00Z" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_vertical_units = "meters" ;
		:geospatial_vertical_positive = "up" ;
		:geospatial_vertical_resolution = 0. ;
		:time_coverage_resolution = "PT1H" ;
		:creator_email = "cheung@hawaii.edu" ;
		:creator_name = "Kwok Fai Cheung" ;
		:creator_url = "http://www.ore.hawaii.edu/OE/cheung_research.htm" ;
		:date_created = "2013-02-19" ;
		:date_issued = "2013-02-19" ;
		:date_modified = "2014-06-23" ;
		:institution = "University of Hawaii" ;
		:project = "Pacific Islands Ocean Observing System (PacIOOS)" ;
		:contributor_name = "Jim Potemra" ;
		:contributor_role = "distributor" ;
		:publisher_email = "info@pacioos.org" ;
		:publisher_name = "Pacific Islands Ocean Observing System (PacIOOS)" ;
		:publisher_url = "http://pacioos.org" ;
		:license = "The data may be used and redistributed for free but is not intended for legal use, since it may contain inaccuracies. Neither the data Contributor, University of Hawaii, PacIOOS, NOAA, State of Hawaii nor the United States Government, nor any of their employees or contractors, makes any warranty, express or implied, including warranties of merchantability and fitness for a particular purpose, or assumes any legal liability for the accuracy, completeness, or usefulness, of this information." ;
		:acknowledgment = "The Pacific Islands Ocean Observing System (PacIOOS) is funded through the National Oceanic and Atmospheric Administration (NOAA) as a Regional Association within the U.S. Integrated Ocean Observing System (IOOS). PacIOOS is coordinated by the University of Hawaii School of Ocean and Earth Science and Technology (SOEST)." ;
		:source = "Simulating WAves Nearshore (SWAN) numerical wave model" ;
		:references = "http://pacioos.org/waves/model-tutuila/, http://swanmodel.sourceforge.net" ;
		:history = "FMRC Best Dataset" ;
}
