
netcdf \3mf07 {
dimensions:
	maxStrlen64 = 64 ;
	profile = 5 ;
	z = 10 ;
variables:
	float latitude(profile) ;
		latitude:long_name = "Profile Location" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:valid_max = "90.0" ;
		latitude:valid_min = "-90.0" ;
		latitude:axis = "Y" ;
		latitude:_CoordinateAxisType = "Lat" ;
		latitude:ioos_category = "Location" ;
		latitude:_FillValue = -9999.9f ;
		latitude:missing_value = -9999.9f ;
	float longitude(profile) ;
		longitude:long_name = "Profile Location" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:valid_max = "180.0" ;
		longitude:valid_min = "-180.0" ;
		longitude:_CoordinateAxisType = "Lon" ;
		longitude:ioos_category = "Location" ;
		longitude:_FillValue = -9999.9f ;
		longitude:missing_value = -9999.9f ;
		longitude:axis = "X" ;
	float z(z) ;
		z:long_name = "Depth" ;
		z:standard_name = "depth" ;
		z:ioos_category = "Location" ;
		z:units = "m" ;
		z:positive = "down" ;
		z:_FillValue = -9999.9f ;
		z:missing_value = -9999.9f ;
		z:coverage_content_type = "physicalMeasurement" ;
		z:comment = "depth was calculated from pressure using Sea-Bird Electronics document AN69, http://www.seabird.com/document/an69-conversion-pressure-depth" ;
		z:axis = "Z" ;
	int flag(profile) ;
		flag:long_name = "flag" ;
		flag:units = "" ;
		flag:missing_value = -9999.9f ;
		flag:coordinates = "time latitude longitude z" ;
	int haul(profile) ;
		haul:long_name = "haul_number" ;
		haul:units = "" ;
		haul:missing_value = -9999.9f ;
		haul:coordinates = "time latitude longitude z" ;
	char file(profile, maxStrlen64) ;
		file:long_name = "file" ;
		file:units = "" ;
		file:missing_value = -9999.9f ;
		file:coordinates = "time latitude longitude z" ;
	int time(profile) ;
		time:long_name = "Profile Time" ;
		time:standard_name = "time" ;
		time:calendar = "standard" ;
		time:units = "seconds since 1970-01-01T00:00:00Z" ;
		time:axis = "T" ;
		time:ioos_category = "Time" ;
		time:time_origin = "01-JAN-1970 00:00:00" ;
		time:_CoordinateAxisType = "Time" ;
		time:missing_value = -9999.9 ;
	char profile(profile, maxStrlen64) ;
		profile:long_name = "Profile Name" ;
		profile:cf_role = "profile_id" ;
	int crs ;
		crs:long_name = "Coordinate Reference System" ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:epsg_code = "4326" ;
		crs:semi_major_axis = "6378137.0" ;
		crs:inverse_flattening = "298.257223563" ;
	float pressure(profile, z) ;
		pressure:long_name = "Sea Water Pressure" ;
		pressure:standard_name = "sea_water_pressure" ;
		pressure:units = "10000.0 Pa" ;
		pressure:_FillValue = -9999.9f ;
		pressure:missing_value = -9999.9f ;
		pressure:coordinates = "time latitude longitude z" ;
		pressure:coverage_content_type = "physicalMeasurement" ;
	float temperature(profile, z) ;
		temperature:long_name = "Water Temperature" ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "degree_Celsius" ;
		temperature:_FillValue = -9999.9f ;
		temperature:missing_value = -9999.9f ;
		temperature:coordinates = "time latitude longitude z" ;
		temperature:coverage_content_type = "physicalMeasurement" ;
	float conductivity(profile, z) ;
		conductivity:long_name = "Conductivity" ;
		conductivity:standard_name = "sea_water_electrical_conductivity" ;
		conductivity:units = "mS.cm-1" ;
		conductivity:_FillValue = -9999.9f ;
		conductivity:missing_value = -9999.9f ;
		conductivity:coordinates = "time latitude longitude z" ;
		conductivity:coverage_content_type = "physicalMeasurement" ;
	float salinity(profile, z) ;
		salinity:long_name = "Salinity" ;
		salinity:standard_name = "sea_water_practical_salinity" ;
		salinity:units = "1e-3" ;
		salinity:_FillValue = -9999.9f ;
		salinity:missing_value = -9999.9f ;
		salinity:coordinates = "time latitude longitude z" ;
		salinity:coverage_content_type = "physicalMeasurement" ;
	float sigma_t(profile, z) ;
		sigma_t:long_name = "Sea Water Sigma Theta" ;
		sigma_t:standard_name = "sea_water_sigma_theta" ;
		sigma_t:units = "kg m-3" ;
		sigma_t:_FillValue = -9999.9f ;
		sigma_t:missing_value = -9999.9f ;
		sigma_t:coordinates = "time latitude longitude z" ;
		sigma_t:comments = "sigma-t is sea water density minus 1000 km m-3" ;
		sigma_t:coverage_content_type = "physicalMeasurement" ;

// global attributes:
		:Conventions = "CF-1.6, ACDD-1.3" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention Standard Name Table v27" ;
		:featureType = "profile" ;
		:cdm_data_type = "Profile" ;
		:nodc_template_version = "NODC_NetCDF_Profile_Incomplete_Template_v1.1" ;
		:cruise = "3MF07" ;
		:platform = "Miller Freeman" ;
		:platform_vocabulary = "" ;
		:vessel_name = "Miller Freeman" ;
		:platform_nodc = "31FN" ;
		:platform_wod = "1544" ;
		:platform_ircs = "WTDM" ;
		:instrument = "Sea-Bird SBE 19" ;
		:instrument_vocabulary = "" ;
		:urn = "urn:ioos:station:gov.noaa.afsc:3mf07" ;
		:id = "3mf07" ;
		:naming_authority = "gov.noaa.afsc" ;
		:data_center_url = "www.pmel.noaa.gov" ;
		:sea_name = "Bering Sea" ;
		:project = "NPCREP" ;
		:title = "3MF07 SeaCAT Data" ;
		:description = "To recover and deploy surface and subsurface oceanographic instrumentation moorings.  To complete Conductivity, Temperature, and Depth (CTD) profiler casts." ;
		:summary = "To recover and deploy surface and subsurface oceanographic instrumentation moorings.  To complete Conductivity, Temperature, and Depth (CTD) profiler casts." ;
		:processing_level = " The raw data are processed using the SeaBird SBE Data Processing software.  The raw data are low pass filtered, aligned to pressure, flagged for wildly incorrect values, averaged to 1 meter bins, and split into up and down casts. Header information about the location and data/time of the cast are added manually.  The upcasts are instpected visually for noisy or erroneous data and those casts are removed." ;
		:keywords = "biological sampling, physical oceanography, salinity, temperature, conductivity, sigma-T, SeaCAT, fish larvae, zooplankton,  mooring deployment, mooring recovery. Utow, Bering Sea, 60cm bongo" ;
		:keywords_vocabulary = "GCMD Earth Science Keywords. Version 5.3.3" ;
		:source = "NOAA/NMFS/AFSC" ;
		:institution = "NOAA/NMFS/AFSC" ;
		:creator_name = "Carol DeWitt" ;
		:creator_url = "www.pmel.noaa.gov" ;
		:creator_email = "" ;
		:creator_institution = "NOAA/NMFS/AFSC" ;
		:netcdf_writer = "Axiom Data Science" ;
		:netcdf_writer_email = "luc@axiomdatascience.com, rob@axiomdatascience.com" ;
		:netcdf_creator_url = "http://www.axiomdatascience.com/" ;
		:netcdf_date_created = "2016-09-13T17:53:49Z" ;
		:date_metadata_modified = "2016-09-13T17:53:49Z" ;
		:date_modified = "" ;
		:references = "" ;
		:date_issued = "2015-12-01T00:00:00Z" ;
		:date_created = "2015-12-01T00:00:00Z" ;
		:contributor_name = "William Floering, Peter Proctor, Steve Smith, Marty Reedy" ;
		:contributor_role = "Scientist" ;
		:publisher_name = "Tiffany C. Vance" ;
		:publisher_institution = "NOAA/NMFS/AFSC" ;
		:publisher_email = "Tiffany.C.Vance@noaa.gov" ;
		:publisher_url = "" ;
		:history = "NetCDF generated by Axiom from excel file provided by Tiffany Vance, NOAA. " ;
		:license = "There are no legal restrictions on access to the data. They reside in public domain and can be freely distributed. User must read and fully comprehend the metadata prior to use. Applications or inferences derived from the data should be carefully considered for accuracy. Data will reside at the Alaska Fisheries Science Center. Acknowledgement of NOAA/NMFS/AFSC, as the source from which these data were obtained in any publications and/or other representations of these, data is suggested." ;
		:metadata_link = "" ;
		:acknowledgment = "Acknowledgement of NOAA/NMFS/AFSC, as the source from which these data were obtained in any publications and/or other representations of these, data is suggested." ;
		:comment = "" ;
		:time_coverage_start = "2007-04-24T15:00:00Z" ;
		:time_coverage_end = "2007-04-24T22:07:00Z" ;
		:time_coverage_duration = 25620000. ;
		:time_coverage_resolution = "point" ;
		:geospatial_bounds = "POLYGON(-163.9 57.8937,-163.023 57.8937,-163.023 57.0008,-163.9 57.0008,-163.9 57.8937)" ;
		:geospatial_bounds_crs = "EPSG:4326" ;
		:geospatial_lat_max = 57.8937 ;
		:geospatial_lat_min = 57.0008 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lat_resolution = "point" ;
		:geospatial_lon_max = -163.023 ;
		:geospatial_lon_min = -163.9 ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lon_resolution = "point" ;
		:geospatial_vertical_positive = "down" ;
		:geospatial_vertical_min = 0.99 ;
		:geospatial_vertical_max = 56.47 ;
		:geospatial_vertical_units = "meters" ;
		:geospatial_vertical_resolution = "1.0" ;
		:geospatial_vertical_reference = "mean_sea_level" ;
		:geospatial_pressure_min = "0.0" ;
		:geospatial_pressure_max = "57.0" ;
		:geospatial_pressure_units = "dbar" ;
		:geospatial_pressure_resolution = "1" ;
}
