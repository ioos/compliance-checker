netcdf index_ragged {
dimensions:
	obs = UNLIMITED ; // (213 currently)
	trajectory = 10 ;
	name_strlen = 50 ;
variables:
	float lat(obs) ;
		lat:units = "degrees_north" ;
		lat:long_name = "station latitude" ;
		lat:standard_name = "latitude" ;
	float lon(obs) ;
		lon:units = "degrees_east" ;
		lon:long_name = "station longitude" ;
		lon:standard_name = "longitude" ;
	int trajectory_info(trajectory) ;
		trajectory_info:long_name = "trajectory info" ;
		trajectory_info:missing_value = -999 ;
	char trajectory_name(trajectory, name_strlen) ;
		trajectory_name:cf_role = "trajectory_id" ;
		trajectory_name:long_name = "trajectory name" ;
	int trajectory_index(obs) ;
		trajectory_index:long_name = "index of trajectory this obs belongs to" ;
		trajectory_index:instance_dimension = "trajectory" ;
	int time(obs) ;
		time:long_name = "time of measurement" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1990-01-01 00:00:00" ;
		time:missing_value = -999 ;
	float z(obs) ;
		z:long_name = "height above mean sea level" ;
		z:standard_name = "altitude" ;
		z:units = "m" ;
		z:positive = "up" ;
		z:axis = "Z" ;
		z:missing_value = -999.9f ;
	float temperature(obs) ;
		temperature:long_name = "Air Temperature" ;
		temperature:standard_name = "air_temperature" ;
		temperature:units = "Celsius" ;
		temperature:coordinates = "time lat lon z" ;
		temperature:missing_value = -999.9f ;
	float humidity(obs) ;
		humidity:long_name = "Humidity" ;
		humidity:standard_name = "specific_humidity" ;
		humidity:units = "Percent" ;
		humidity:coordinates = "time lat lon z" ;
		humidity:missing_value = -999.9f ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:featureType = "trajectory" ;
data:

 lat = 11.25615, 26.10413, 22.41421, 22.18116, 2.177301, 14.65077, 8.425178,
    33.27557, 7.699538, 12.65807, 22.59023, 35.84382, 41.75186, 44.95267,
    41.49166, 31.4028, 20.86521, 29.92925, 40.79485, 7.187255, 37.35788,
    17.61622, 29.03985, 44.19264, 21.68499, 22.39728, 12.24242, 26.04828,
    29.84989, 11.87822, 0.4776838, 35.66367, 31.27619, 23.92727, 12.09872,
    3.706677, 13.97815, 2.305441, 0.1856368, 0.3515074, 36.93685, 25.41243,
    30.47535, 17.78078, 7.249343, 24.00756, 44.45137, 36.97704, 30.41355,
    39.9559, 7.445425, 21.05626, 5.065194, 2.547434, 3.349946, 23.44335,
    2.681866, 18.70734, 4.612935, 2.512696, 37.66089, 30.70432, 42.76654,
    33.08486, 6.084778, 39.70843, 28.33197, 1.223405, 38.01586, 3.699682,
    2.316901, 35.92374, 30.71458, 20.204, 4.404234, 13.65772, 22.67983,
    17.34453, 15.95195, 19.13686, 43.36827, 36.43596, 16.88155, 5.257358,
    7.246674, 1.400879, 15.63431, 42.32153, 15.68266, 33.21914, 40.09315,
    28.85555, 20.94757, 12.3212, 36.19291, 30.34604, 32.3859, 30.51254,
    3.334529, 11.59718, 8.42951, 28.87055, 3.602655, 34.14508, 37.11425,
    41.03566, 24.49625, 6.173713, 8.171118, 32.33793, 37.4291, 24.66317,
    40.02692, 40.21726, 2.723573, 27.94735, 28.4283, 20.29399, 33.83424,
    33.06853, 21.15303, 12.59542, 37.33821, 37.76236, 30.25255, 13.93048,
    1.547064, 7.328507, 9.377513, 29.12751, 3.766602, 40.7905, 16.42247,
    35.71611, 15.67354, 26.41485, 8.666093, 3.303721, 3.405675, 19.47607,
    20.71446, 9.468412, 36.72459, 3.348803, 44.85631, 39.74762, 29.31821,
    4.541548, 11.51457, 41.51421, 40.40759, 4.126002, 36.88403, 22.56794,
    16.48313, 38.77134, 32.14177, 17.71075, 3.117972, 2.657588, 15.24631,
    2.316706, 9.206306, 6.183945, 19.74638, 3.791813, 32.1823, 0.7473986,
    34.80326, 2.932063, 24.79398, 31.73436, 10.17321, 44.13942, 0.4635795,
    32.58381, 2.969093, 0.7101297, 6.049965, 23.23353, 19.27657, 37.33231,
    6.420473, 24.66804, 0.8633785, 42.47254, 43.24734, 25.53198, 43.51039,
    10.20917, 30.8017, 21.22977, 15.69756, 20.59331, 31.61997, 16.75511,
    5.537777, 44.28425, 22.34849, 6.084063, 36.75227, 13.18288, 25.23589,
    42.4052, 8.214571, 15.91778, 40.54069, 1.812273, 21.60521, 41.05975,
    26.5076, 19.88841, 38.60466 ;

 lon = -5.989336, -2.662698, -23.53803, -34.35585, -58.38861, -52.61451,
    -0.7129942, -52.05439, -34.31932, -42.76257, -15.92119, -46.72515,
    -44.9617, -63.97917, -41.69743, -8.890802, -31.29523, -61.6931,
    -52.59704, -50.17197, -37.69957, -57.86943, -70.20708, -58.25657,
    -46.1655, -53.94893, -75.69691, -8.550176, -38.24889, -3.490612,
    -39.24084, -3.612438, -47.12128, -48.02716, -55.01497, -59.63803,
    -38.12038, -50.87202, -30.13649, -14.03829, -7.792219, -72.6375,
    -20.88588, -53.71122, -55.1488, -41.42715, -1.574568, -37.43023,
    -7.373155, -29.56204, -50.04349, -20.28753, -36.01645, -7.64748,
    -49.57981, -2.64897, -9.46538, -46.31868, -2.049518, -64.91229,
    -68.88179, -42.89665, -51.48783, -6.27085, -62.04066, -30.79151,
    -2.580461, -21.22981, -7.61332, -16.17166, -23.74372, -61.22404,
    -72.97459, -20.26349, -20.53997, -3.180203, -49.06118, -37.38556,
    -65.62891, -13.13425, -67.3617, -62.12461, -15.67471, -15.32692,
    -40.40166, -72.79348, -28.02558, -31.81828, -1.080388, -67.15468,
    -72.98028, -17.48965, -61.34195, -35.70835, -1.923249, -21.76571,
    -12.04998, -74.69545, -30.8238, -75.83024, -57.93318, -30.22355,
    -71.86282, -34.07526, -18.59933, -52.08774, -6.3491, -52.88477,
    -15.02928, -41.72115, -10.90716, -13.49223, -66.11868, -19.19154,
    -24.1513, -28.1119, -33.80967, -23.85966, -69.89976, -59.48049, -57.7855,
    -56.86527, -45.3292, -21.1472, -20.11768, -32.99857, -26.61098,
    -34.56091, -58.16519, -65.28774, -3.262689, -27.42458, -44.577,
    -18.71307, -75.23668, -50.39792, -37.36423, -59.43841, -13.20477,
    -43.58611, -8.478054, -19.66856, -14.8859, -31.48991, -62.27028,
    -61.14234, -53.99629, -58.88906, -31.54302, -35.90159, -54.26013,
    -41.56313, -59.35286, -49.54479, -57.84679, -2.264266, -7.235641,
    -64.94084, -65.73678, -54.36418, -64.24323, -52.50892, -71.1492,
    -4.25458, -10.47351, -37.3678, -69.27312, -29.40901, -16.01023,
    -12.14635, -41.12995, -56.01423, -65.60724, -74.3843, -69.52895,
    -69.94255, -46.57818, -6.044638, -73.67628, -36.0216, -47.81919,
    -46.84343, -21.60306, -7.668083, -68.5562, -70.67887, -34.45117,
    -60.26342, -64.72975, -40.86289, -26.85923, -61.6675, -52.7378,
    -72.34982, -7.364043, -18.06771, -34.36699, -65.99042, -52.3617,
    -45.11955, -74.25336, -40.7113, -41.43104, -30.44535, -18.81168,
    -26.02182, -15.331, -29.46848, -58.86243, -63.42926, -10.08484,
    -26.79434, -1.817341 ;

 trajectory_info = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9 ;

 trajectory_name =
  "Trajectory0",
  "Trajectory1",
  "Trajectory2",
  "Trajectory3",
  "Trajectory4",
  "Trajectory5",
  "Trajectory6",
  "Trajectory7",
  "Trajectory8",
  "Trajectory9" ;

 trajectory_index = 8, 3, 4, 4, 5, 4, 7, 2, 9, 0, 3, 4, 1, 7, 9, 3, 3, 4, 9,
    9, 9, 7, 9, 8, 3, 4, 7, 3, 9, 0, 4, 2, 6, 3, 1, 8, 4, 2, 8, 9, 5, 4, 7,
    0, 0, 0, 7, 0, 2, 7, 7, 3, 1, 0, 6, 1, 2, 1, 0, 9, 6, 1, 6, 5, 2, 3, 4,
    9, 2, 9, 1, 9, 0, 7, 6, 3, 4, 8, 2, 9, 3, 7, 8, 6, 7, 6, 7, 5, 1, 1, 3,
    3, 7, 1, 3, 0, 9, 2, 7, 6, 8, 1, 1, 4, 1, 9, 7, 4, 2, 9, 6, 0, 4, 7, 0,
    7, 7, 3, 1, 7, 1, 7, 4, 9, 9, 6, 5, 6, 4, 8, 9, 7, 0, 5, 7, 9, 5, 8, 4,
    1, 2, 9, 8, 0, 7, 2, 4, 0, 3, 5, 2, 0, 6, 4, 7, 4, 6, 0, 4, 4, 6, 7, 2,
    8, 6, 6, 4, 2, 1, 7, 7, 1, 3, 2, 7, 9, 8, 4, 2, 1, 2, 7, 1, 7, 2, 1, 5,
    6, 7, 8, 5, 8, 9, 8, 9, 2, 3, 3, 3, 5, 7, 6, 9, 2, 1, 9, 2, 5, 0, 1, 9,
    5, 0 ;

 time = 72000, 111600, 68400, 122400, 162000, 144000, 57600, 36000, 68400,
    118800, 21600, 43200, 28800, 108000, 154800, 10800, 136800, 158400,
    46800, 158400, 104400, 176400, 36000, 104400, 82800, 28800, 158400,
    118800, 133200, 136800, 64800, 79200, 90000, 50400, 90000, 144000, 18000,
    36000, 122400, 165600, 172800, 169200, 86400, 3600, 118800, 129600,
    115200, 100800, 25200, 129600, 108000, 64800, 21600, 10800, 21600, 18000,
    36000, 169200, 79200, 68400, 158400, 54000, 28800, 64800, 46800, 147600,
    169200, 111600, 79200, 100800, 151200, 154800, 39600, 126000, 46800,
    25200, 136800, 7200, 97200, 79200, 165600, 162000, 118800, 0, 25200,
    169200, 169200, 72000, 133200, 122400, 154800, 169200, 82800, 18000,
    133200, 144000, 64800, 104400, 68400, 72000, 154800, 90000, 75600, 10800,
    32400, 97200, 46800, 172800, 90000, 133200, 3600, 25200, 151200, 36000,
    75600, 129600, 151200, 108000, 111600, 151200, 172800, 3600, 28800,
    68400, 136800, 90000, 93600, 0, 176400, 82800, 86400, 165600, 154800,
    39600, 93600, 115200, 21600, 43200, 61200, 93600, 61200, 50400, 104400,
    158400, 147600, 75600, 0, 133200, 0, 126000, 50400, 140400, 108000,
    147600, 25200, 126000, 90000, 165600, 100800, 86400, 3600, 97200, 72000,
    118800, 144000, 54000, 21600, 86400, 162000, 86400, 154800, 122400,
    28800, 93600, 28800, 43200, 172800, 18000, 165600, 151200, 3600, 25200,
    54000, 162000, 133200, 28800, 18000, 43200, 86400, 176400, 172800,
    104400, 18000, 14400, 151200, 36000, 111600, 3600, 133200, 154800,
    147600, 50400, 0, 158400, 118800, 176400, 133200, 133200, 154800, 129600,
    136800, 86400, 14400 ;

 z = 12.51808, 7.372036, 5.799932, 20.12702, 1.764841, 19.18218, 4.44464,
    0.03310063, 29.50963, 8.532058, 16.35266, 13.58115, 28.27637, 4.366767,
    20.38323, 3.586328, 11.11897, 22.30022, 16.46136, 16.86729, 4.325697,
    16.50045, 2.312687, 25.4671, 26.26118, 22.33489, 29.15273, 17.85277,
    13.19439, 5.735756, 22.62788, 9.360034, 12.95132, 11.07303, 7.477769,
    28.16613, 27.99436, 22.90513, 28.66971, 15.94959, 21.66013, 14.11007,
    25.57854, 16.84065, 0.415791, 12.5649, 2.325282, 1.742066, 24.94547,
    16.64068, 26.13454, 13.14445, 8.728339, 20.30043, 20.88193, 0.08922961,
    11.32374, 19.46538, 23.49089, 23.33969, 16.94271, 13.68294, 28.23238,
    5.902096, 13.79568, 0.3863254, 16.6489, 7.460392, 1.204016, 21.68154,
    17.06803, 12.06111, 15.4019, 26.2678, 9.876749, 29.56433, 14.53347,
    6.870228, 29.69398, 2.245085, 28.9268, 4.583749, 29.69282, 13.04906,
    1.512483, 22.88785, 13.26198, 22.86892, 12.05387, 21.77244, 20.18067,
    20.21082, 18.28759, 9.992888, 4.024284, 11.44874, 18.03653, 0.142246,
    24.32986, 21.6673, 22.37223, 24.45863, 1.028929, 11.27909, 12.96912,
    29.51361, 16.17835, 16.55074, 16.81288, 0.9152418, 4.687667, 12.44715,
    15.05259, 23.95142, 8.311193, 5.329725, 9.22603, 2.188019, 5.634934,
    14.02315, 2.931201, 21.93977, 8.667504, 21.51781, 0.1166571, 8.247705,
    15.02659, 17.7737, 0.7352603, 5.177349, 24.14933, 15.98668, 6.480564,
    5.164011, 9.530041, 21.05122, 18.45421, 7.870076, 0.4085527, 8.535103,
    17.55896, 16.71356, 10.36592, 10.28535, 10.61128, 7.40977, 0.4369197,
    8.551613, 20.86436, 2.689621, 23.69171, 24.28577, 26.60997, 9.152925,
    5.37336, 10.43244, 29.37995, 0.6106723, 24.26659, 23.86881, 21.48618,
    0.09007654, 18.17645, 4.797531, 7.067278, 14.12353, 13.73014, 27.95491,
    3.776026, 16.52352, 1.692304, 11.92638, 25.06545, 10.02483, 28.19705,
    9.880977, 3.647643, 1.075158, 19.46502, 3.479654, 24.82868, 26.67636,
    24.10556, 7.428996, 28.01834, 10.31546, 11.68204, 23.85533, 28.76868,
    9.559212, 6.03133, 2.056599, 12.88738, 14.75593, 13.85003, 25.33521,
    23.70653, 24.96098, 24.8398, 17.94507, 6.896889, 17.03668, 28.3191,
    29.14639, 7.3838, 4.964994, 9.436576, 21.62823, 20.98346, 11.14172,
    7.991476, 29.63633, 22.9028 ;

 temperature = 14.90271, 24.24385, 1.494066, 6.831084, 27.893, 33.67621,
    20.69297, 19.61122, 17.45888, 1.446625, 5.125631, 35.8677, 12.99567,
    28.21161, 31.1266, 12.29142, 39.75038, 6.404823, 17.65268, 23.69756,
    14.05361, 13.79113, 29.22715, 24.8389, 22.293, 18.33682, 34.71552,
    21.25107, 27.40752, 19.85405, 1.102716, 26.13454, 20.0989, 34.58173,
    10.09682, 34.69993, 21.41687, 24.60953, 2.707067, 28.78928, 36.26309,
    7.720104, 20.29351, 6.168052, 16.10084, 37.99405, 0.5267054, 15.17727,
    16.9081, 2.68189, 21.16533, 35.04569, 8.063735, 16.21928, 4.422824,
    7.724518, 17.27993, 39.00298, 32.56659, 14.87465, 15.83106, 13.7587,
    13.87703, 38.87086, 3.104527, 27.18122, 3.531546, 38.92941, 32.89718,
    15.72652, 9.8498, 30.11894, 35.62276, 6.708208, 32.10239, 15.3041,
    25.26304, 34.48993, 20.19512, 0.2903271, 3.622684, 2.85062, 12.61744,
    23.07567, 0.5586658, 22.41853, 22.86525, 3.229707, 3.379141, 8.767585,
    9.436486, 9.661129, 33.93568, 28.27926, 28.42878, 23.78411, 17.47237,
    29.69628, 7.52533, 3.482231, 6.826304, 21.11233, 2.944838, 36.02184,
    16.79605, 13.76455, 38.61915, 33.59118, 20.93422, 16.73082, 37.01011,
    9.472145, 0.05421121, 35.55663, 14.59343, 17.78524, 10.66914, 31.76535,
    22.87287, 15.78297, 30.92633, 1.031407, 32.86114, 19.20944, 35.08533,
    14.45549, 5.093784, 4.045129, 36.97565, 16.91204, 25.10888, 1.929165,
    36.06869, 16.66244, 31.84952, 3.524928, 1.354704, 10.48365, 27.1373,
    12.30132, 2.691948, 27.47651, 13.98832, 16.22222, 4.994209, 31.78442,
    13.77028, 2.929394, 29.53318, 31.14371, 11.47821, 31.36297, 22.94642,
    24.2277, 16.57454, 32.16871, 19.67619, 5.641278, 3.958635, 31.70868,
    30.52293, 20.18705, 39.97938, 30.04643, 17.13696, 3.175597, 1.988845,
    27.89935, 32.00631, 16.65858, 18.483, 9.31581, 19.38959, 39.51171,
    24.08715, 16.227, 22.69785, 36.4146, 1.840191, 11.65769, 36.54749,
    12.34812, 37.90659, 28.72273, 12.70363, 34.74529, 12.26348, 2.720131,
    2.401074, 6.551149, 25.93415, 29.62659, 21.72955, 16.11036, 2.032868,
    1.986544, 14.58139, 10.11439, 10.15086, 22.30464, 17.00665, 39.1347,
    21.63502, 3.290949, 38.27164, 21.9019, 17.38786, 22.71373, 25.47452,
    32.77483, 38.94097, 21.50251, 23.38549 ;

 humidity = 37.23755, 12.86247, 20.66832, 55.93755, 28.2276, 47.91003,
    46.91182, 70.05315, 64.52536, 35.24868, 6.144204, 25.3432, 35.19174,
    6.857599, 73.46922, 68.64112, 31.69522, 16.41469, 32.78758, 44.50916,
    19.58626, 67.18636, 38.4418, 29.44308, 58.00679, 21.86452, 51.05852,
    45.4691, 8.350641, 18.38804, 44.15499, 64.43467, 64.32681, 19.34761,
    0.09478192, 62.03254, 21.54085, 52.27968, 32.77289, 68.97393, 20.62231,
    20.59801, 65.2218, 79.25449, 69.70883, 54.40137, 15.02394, 17.44944,
    61.93802, 71.51801, 11.04534, 7.114886, 10.6127, 15.91914, 1.093509,
    40.47393, 31.31579, 61.54602, 32.63131, 58.71174, 74.66438, 29.86826,
    44.8269, 6.804867, 51.10857, 47.32163, 39.24802, 29.47629, 49.44198,
    12.47171, 54.50966, 66.37208, 79.22325, 73.69112, 59.76095, 28.07529,
    40.53505, 61.64103, 1.367835, 29.19541, 24.63598, 13.36296, 19.15088,
    17.24242, 58.86948, 10.36386, 15.20454, 56.35379, 8.099169, 23.769,
    24.79614, 14.69656, 50.11193, 25.35903, 59.18938, 51.97684, 44.87966,
    56.51338, 76.7057, 37.08824, 18.17326, 36.34776, 57.81669, 15.94002,
    31.54479, 66.87031, 12.56461, 67.00338, 58.19665, 57.84406, 22.33975,
    51.16273, 16.50468, 11.02816, 79.05337, 68.78816, 37.46039, 31.49598,
    66.92045, 53.46638, 35.19886, 49.43015, 29.39922, 13.55865, 71.05666,
    13.83892, 45.22563, 0.02646556, 15.81763, 63.98837, 0.5120609, 10.33802,
    53.50613, 24.63119, 6.965268, 47.22089, 36.78447, 35.98283, 35.40593,
    34.8849, 49.4609, 53.93727, 3.188482, 66.85195, 44.25605, 45.74578,
    45.21314, 39.30257, 0.7206169, 54.77544, 22.18368, 51.29797, 38.16368,
    73.97604, 35.80253, 71.73385, 50.23185, 9.621942, 74.90228, 78.32967,
    8.03379, 10.05789, 79.54096, 38.2582, 26.61588, 36.16071, 7.350058,
    25.95598, 14.06559, 75.5065, 65.43004, 78.54383, 48.77426, 18.51248,
    71.97946, 45.68407, 26.03132, 51.98213, 23.95672, 74.53979, 43.14886,
    49.58644, 27.06123, 25.66633, 28.73472, 60.32231, 49.05508, 16.17089,
    11.29831, 24.5825, 15.77298, 0.8424936, 13.64856, 55.91599, 38.14489,
    44.76837, 68.57007, 2.255769, 50.99001, 30.59435, 36.69022, 25.05376,
    28.26003, 10.82617, 5.319588, 22.8674, 38.64904, 67.63327, 63.17289,
    66.06119, 69.17253, 18.88459, 10.31085 ;
}
