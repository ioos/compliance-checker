netcdf temp {
dimensions:
	TIME = UNLIMITED ; // (22 currently)
	h_num = 15 ;
	h_string = 236 ;
variables:
	double TIME(TIME) ;
		TIME:standard_name = "time" ;
		TIME:long_name = "time" ;
		TIME:units = "days since 1950-01-01 00:00:00Z" ;
		TIME:axis = "T" ;
		TIME:valid_min = 0. ;
		TIME:valid_max = 90000. ;
		TIME:_FillValue = -9999. ;
		TIME:comment = "Relative julian days with decimal part as parts \n",
			"of the day" ;
		TIME:calendar = "gregorian" ;
	float LATITUDE(TIME) ;
		LATITUDE:standard_name = "latitude" ;
		LATITUDE:long_name = "latitude" ;
		LATITUDE:units = "degrees_north" ;
		LATITUDE:axis = "Y" ;
		LATITUDE:valid_min = -90.f ;
		LATITUDE:valid_max = 90.f ;
		LATITUDE:_FillValue = -9999.f ;
		LATITUDE:reference_datum = "geographical coordinates, WGS84" ;
		LATITUDE:coordinates = "TIME LATITUDE LONGITUDE" ;
	float LONGITUDE(TIME) ;
		LONGITUDE:standard_name = "longitude" ;
		LONGITUDE:long_name = "longitude" ;
		LONGITUDE:units = "degrees_east" ;
		LONGITUDE:axis = "X" ;
		LONGITUDE:valid_min = -180.f ;
		LONGITUDE:valid_max = 180.f ;
		LONGITUDE:_FillValue = -9999.f ;
		LONGITUDE:reference_datum = "geographical coordinates, WGS84" ;
		LONGITUDE:coordinates = "TIME LATITUDE LONGITUDE" ;
	float PL_CMP(TIME) ;
		PL_CMP:long_name = "compass direction" ;
		PL_CMP:units = "degrees_north" ;
		PL_CMP:observation_type = "measured" ;
		PL_CMP:_FillValue = -9999.f ;
		PL_CMP:coordinates = "TIME LATITUDE LONGITUDE" ;
	float PL_CRS(TIME) ;
		PL_CRS:standard_name = "platform_course" ;
		PL_CRS:long_name = "platform course" ;
		PL_CRS:units = "degree" ;
		PL_CRS:observation_type = "measured" ;
		PL_CRS:_FillValue = -9999.f ;
		PL_CRS:comment = "(clockwise from true north)" ;
		PL_CRS:coordinates = "TIME LATITUDE LONGITUDE" ;
	float PL_SPD(TIME) ;
		PL_SPD:standard_name = "platform_speed_wrt_ground" ;
		PL_SPD:long_name = "platform speed over ground" ;
		PL_SPD:units = "meter second-1" ;
		PL_SPD:observation_type = "measured" ;
		PL_SPD:_FillValue = -9999.f ;
		PL_SPD:coordinates = "TIME LATITUDE LONGITUDE" ;
	float WDIR(TIME) ;
		WDIR:standard_name = "wind_to_direction" ;
		WDIR:long_name = "earth relative wind direction (oceanographic)" ;
		WDIR:units = "degree" ;
		WDIR:_FillValue = -9999.f ;
		WDIR:observation_type = "calculated" ;
		WDIR:coordinates = "TIME LATITUDE LONGITUDE" ;
	float WSPD(TIME) ;
		WSPD:standard_name = "wind_speed" ;
		WSPD:long_name = "earth relative wind speed" ;
		WSPD:units = "meter second-1" ;
		WSPD:_FillValue = -9999.f ;
		WSPD:observation_type = "calculated" ;
		WSPD:ancillary_variables = "WIND_FLAG" ;
		WSPD:coordinates = "TIME LATITUDE LONGITUDE" ;
	float WIND_H(TIME) ;
		WIND_H:long_name = "wind measurement height above water level" ;
		WIND_H:units = "meter" ;
		WIND_H:_FillValue = -9999.f ;
		WIND_H:coordinates = "TIME LATITUDE LONGITUDE" ;
	short WIND_FLAG(TIME) ;
		WIND_FLAG:long_name = "wind sensor flag" ;
		WIND_FLAG:comment = "1 - mainmast sensor" ;
		WIND_FLAG:flag_meanings = "mainmast_sensor" ;
		WIND_FLAG:flag_values = "1" ;
		WIND_FLAG:coordinates = "TIME LATITUDE LONGITUDE" ;
	float ATMP(TIME) ;
		ATMP:standard_name = "air_pressure" ;
		ATMP:long_name = "atmospheric pressure" ;
		ATMP:units = "hectopascal" ;
		ATMP:_FillValue = -9999.f ;
		ATMP:mslp_indicator = "adjusted to sea level" ;
		ATMP:observation_type = "measured" ;
		ATMP:ancillary_variables = "ATMP_FLAG" ;
		ATMP:coordinates = "TIME LATITUDE LONGITUDE" ;
	float ATMP_H(TIME) ;
		ATMP_H:long_name = "atmospheric pressure measurement height above water level" ;
		ATMP_H:units = "meter" ;
		ATMP_H:_FillValue = -9999.f ;
		ATMP_H:coordinates = "TIME LATITUDE LONGITUDE" ;
	short ATMP_FLAG(TIME) ;
		ATMP_FLAG:long_name = "air pressure sensor flag" ;
		ATMP_FLAG:comment = "1 - currently available the only sensor" ;
		ATMP_FLAG:flag_meanings = "currently_available_the_only_sensor" ;
		ATMP_FLAG:flag_values = 1b ;
		ATMP_FLAG:coordinates = "TIME LATITUDE LONGITUDE" ;
	float AIRT(TIME) ;
		AIRT:standard_name = "air_temperature" ;
		AIRT:long_name = "air temperature" ;
		AIRT:units = "celsius" ;
		AIRT:_FillValue = -9999.f ;
		AIRT:observation_type = "measured" ;
		AIRT:ancillary_variables = "AIRT_FLAG" ;
		AIRT:coordinates = "TIME LATITUDE LONGITUDE" ;
	float AIRT_H(TIME) ;
		AIRT_H:long_name = "air temperature measurement height above water level" ;
		AIRT_H:units = "meter" ;
		AIRT_H:coordinates = "TIME LATITUDE LONGITUDE" ;
	short AIRT_FLAG(TIME) ;
		AIRT_FLAG:long_name = "air temperature sensor flag" ;
		AIRT_FLAG:comment = "1 - currently available the only sensor" ;
		AIRT_FLAG:flag_meanings = "currently_available_the_only_sensor" ;
		AIRT_FLAG:flag_values = 1b ;
		AIRT_FLAG:coordinates = "TIME LATITUDE LONGITUDE" ;
	float RELH(TIME) ;
		RELH:standard_name = "relative_humidity" ;
		RELH:long_name = "relative humidity " ;
		RELH:units = "percent" ;
		RELH:_FillValue = -9999.f ;
		RELH:observation_type = "measured" ;
		RELH:ancillary_variables = "RELH_FLAG" ;
		RELH:coordinates = "TIME LATITUDE LONGITUDE" ;
	float RELH_H(TIME) ;
		RELH_H:long_name = "relative humidity measurement height above water level" ;
		RELH_H:units = "meter" ;
		RELH_H:_FillValue = -9999.f ;
		RELH_H:coordinates = "TIME LATITUDE LONGITUDE" ;
	short RELH_FLAG(TIME) ;
		RELH_FLAG:long_name = "relative humidity sensor flag" ;
		RELH_FLAG:comment = "1 - currently available the only sensor" ;
		RELH_FLAG:flag_meanings = "currently_available_the_only_sensor" ;
		RELH_FLAG:flag_values = 1b ;
		RELH_FLAG:coordinates = "TIME LATITUDE LONGITUDE" ;
	float TEMP(TIME) ;
		TEMP:standard_name = "sea_water_temperature" ;
		TEMP:long_name = "sea water temperature from TSG" ;
		TEMP:units = "celsius" ;
		TEMP:_FillValue = -9999.f ;
		TEMP:observation_type = "measured" ;
		TEMP:ancillary_variables = "TEMP_FLAG" ;
		TEMP:coordinates = "TIME LATITUDE LONGITUDE" ;
	float TEMP_H(TIME) ;
		TEMP_H:long_name = "sea water temeperature measurement depth" ;
		TEMP_H:units = "meter" ;
		TEMP_H:_FillValue = -9999.f ;
		TEMP_H:coordinates = "TIME LATITUDE LONGITUDE" ;
	short TEMP_FLAG(TIME) ;
		TEMP_FLAG:long_name = "sea water temeperature sensor flag" ;
		TEMP_FLAG:comment = "1 - currently available the only sensor" ;
		TEMP_FLAG:flag_meanings = "currently_available_the_only_sensor" ;
		TEMP_FLAG:flag_values = 1b ;
		TEMP_FLAG:coordinates = "TIME LATITUDE LONGITUDE" ;
	float RAIN_AMOUNT(TIME) ;
		RAIN_AMOUNT:standard_name = "rainfall_rate" ;
		RAIN_AMOUNT:long_name = "rain rate" ;
		RAIN_AMOUNT:units = "millimeters hour-1" ;
		RAIN_AMOUNT:_FillValue = -9999.f ;
		RAIN_AMOUNT:observation_type = "measured" ;
		RAIN_AMOUNT:ancillary_variables = "RAIN_AMOUNT_FLAG" ;
		RAIN_AMOUNT:coordinates = "TIME LATITUDE LONGITUDE" ;
	float RAIN_AMOUNT_H(TIME) ;
		RAIN_AMOUNT_H:long_name = "precipitation measurement height above water level" ;
		RAIN_AMOUNT_H:units = "meter" ;
		RAIN_AMOUNT_H:_FillValue = -9999.f ;
		RAIN_AMOUNT_H:coordinates = "TIME LATITUDE LONGITUDE" ;
	short RAIN_AMOUNT_FLAG(TIME) ;
		RAIN_AMOUNT_FLAG:long_name = "precipitation sensor flag" ;
		RAIN_AMOUNT_FLAG:comment = "1 - currently available the only sensor" ;
		RAIN_AMOUNT_FLAG:flag_meanings = "currently_available_the_only_sensor" ;
		RAIN_AMOUNT_FLAG:flag_values = 1b ;
		RAIN_AMOUNT_FLAG:coordinates = "TIME LATITUDE LONGITUDE" ;
	float SW(TIME) ;
		SW:standard_name = "surface_downwelling_shortwave_flux_in_air" ;
		SW:long_name = "short wave radiation" ;
		SW:units = "watts meter-2" ;
		SW:_FillValue = -9999.f ;
		SW:observation_type = "measured" ;
		SW:ancillary_variables = "SW_FLAG" ;
		SW:coordinates = "TIME LATITUDE LONGITUDE" ;
	float SW_H(TIME) ;
		SW_H:long_name = "short-wave radiation measurement height above water level" ;
		SW_H:units = "meter" ;
		SW_H:_FillValue = -9999.f ;
		SW_H:coordinates = "TIME LATITUDE LONGITUDE" ;
	short SW_FLAG(TIME) ;
		SW_FLAG:long_name = "short-wave radiation sensor flag" ;
		SW_FLAG:comment = "1 - starboard sensor, 2 - port sensor" ;
		SW_FLAG:flag_meanings = "starboard_sensor port_sensor" ;
		SW_FLAG:flag_values = 1b, 2b ;
		SW_FLAG:coordinates = "TIME LATITUDE LONGITUDE" ;
	float LW(TIME) ;
		LW:standard_name = "surface_downwelling_longwave_flux_in_air" ;
		LW:long_name = "long wave radiation" ;
		LW:units = "watts meter-2" ;
		LW:_FillValue = -9999.f ;
		LW:observation_type = "measured" ;
		LW:ancillary_variables = "LW_FLAG" ;
		LW:coordinates = "TIME LATITUDE LONGITUDE" ;
	float LW_H(TIME) ;
		LW_H:long_name = "long-wave radiation measurement height above water level" ;
		LW_H:units = "meter" ;
		LW_H:_FillValue = -9999.f ;
		LW_H:coordinates = "TIME LATITUDE LONGITUDE" ;
	byte LW_FLAG(TIME) ;
		LW_FLAG:long_name = "long-wave radiation sensor flag" ;
		LW_FLAG:comment = "1 - starboard sensor, 2 - port sensor, 3 - average of both sensors" ;
		LW_FLAG:flag_meanings = "starboard_sensor port_sensor average_of_both_sensors" ;
		LW_FLAG:flag_values = 1b, 2b, 3b ;
		LW_FLAG:coordinates = "TIME LATITUDE LONGITUDE" ;
	float HS(TIME) ;
		HS:standard_name = "surface_upward_sensible_heat_flux" ;
		HS:long_name = "sensible heat flux" ;
		HS:units = "watts meter-2" ;
		HS:_FillValue = -9999.f ;
		HS:observation_type = "calculated" ;
		HS:coordinates = "TIME LATITUDE LONGITUDE" ;
	float HL(TIME) ;
		HL:standard_name = "surface_upward_latent_heat_flux" ;
		HL:long_name = "latent heat flux" ;
		HL:units = "watts meter-2" ;
		HL:_FillValue = -9999.f ;
		HL:observation_type = "calculated" ;
		HL:coordinates = "TIME LATITUDE LONGITUDE" ;
	float H_RAIN(TIME) ;
		H_RAIN:long_name = "upward heat flux due to rainfall" ;
		H_RAIN:units = "watts meter-2" ;
		H_RAIN:_FillValue = -9999.f ;
		H_RAIN:observation_type = "calculated" ;
		H_RAIN:coordinates = "TIME LATITUDE LONGITUDE" ;
	float TAU(TIME) ;
		TAU:standard_name = "magnitude_of_surface_downward_stress" ;
		TAU:long_name = "wind stress" ;
		TAU:units = "pascal" ;
		TAU:_FillValue = -9999.f ;
		TAU:observation_type = "calculated" ;
		TAU:coordinates = "TIME LATITUDE LONGITUDE" ;
	float SST(TIME) ;
		SST:standard_name = "sea_surface_skin_temperature" ;
		SST:long_name = "sea skin temperature" ;
		SST:units = "celsius" ;
		SST:_FillValue = -9999.f ;
		SST:observation_type = "calculated" ;
		SST:coordinates = "TIME LATITUDE LONGITUDE" ;
	float HEAT_NET(TIME) ;
		HEAT_NET:standard_name = "upward_heat_flux_in_air" ;
		HEAT_NET:long_name = "net heat flux" ;
		HEAT_NET:units = "watts meter-2" ;
		HEAT_NET:_FillValue = -9999.f ;
		HEAT_NET:observation_type = "calculated" ;
		HEAT_NET:coordinates = "TIME LATITUDE LONGITUDE" ;
	float MASS_NET(TIME) ;
		MASS_NET:standard_name = "upward_mass_flux_of_air" ;
		MASS_NET:long_name = "net mass flux" ;
		MASS_NET:units = "kilogram meter-2 second-1" ;
		MASS_NET:_FillValue = -9999.f ;
		MASS_NET:observation_type = "calculated" ;
		MASS_NET:coordinates = "TIME LATITUDE LONGITUDE" ;
	float LW_NET(TIME) ;
		LW_NET:standard_name = "surface_net_upward_longwave_flux" ;
		LW_NET:long_name = "net long-wave radiation" ;
		LW_NET:units = "watts meter-2" ;
		LW_NET:_FillValue = -9999.f ;
		LW_NET:observation_type = "calculated" ;
		LW_NET:coordinates = "TIME LATITUDE LONGITUDE" ;
	float SW_NET(TIME) ;
		SW_NET:standard_name = "surface_net_upward_shortwave_flux" ;
		SW_NET:long_name = "net short-wave radiation" ;
		SW_NET:units = "watts meter-2" ;
		SW_NET:_FillValue = -9999.f ;
		SW_NET:observation_type = "calculated" ;
		SW_NET:coordinates = "TIME LATITUDE LONGITUDE" ;
	float WSPD10M(TIME) ;
		WSPD10M:standard_name = "wind_speed" ;
		WSPD10M:long_name = "calculated neutral wind speed at 10 meters" ;
		WSPD10M:units = "meter second-1" ;
		WSPD10M:_FillValue = -9999.f ;
		WSPD10M:observation_type = "calculated" ;
		WSPD10M:coordinates = "TIME LATITUDE LONGITUDE" ;
	float AIRT1_5M(TIME) ;
		AIRT1_5M:standard_name = "air_temperature" ;
		AIRT1_5M:long_name = "calculated air temperature at 1.5 meters" ;
		AIRT1_5M:units = "celsius" ;
		AIRT1_5M:_FillValue = -9999.f ;
		AIRT1_5M:observation_type = "calculated" ;
		AIRT1_5M:coordinates = "TIME LATITUDE LONGITUDE" ;
	float AIRT2_0M(TIME) ;
		AIRT2_0M:standard_name = "air_temperature" ;
		AIRT2_0M:long_name = "calculated air temperature at 2.0 meters" ;
		AIRT2_0M:units = "celsius" ;
		AIRT2_0M:_FillValue = -9999.f ;
		AIRT2_0M:observation_type = "calculated" ;
		AIRT2_0M:coordinates = "TIME LATITUDE LONGITUDE" ;
	float RELH1_5M(TIME) ;
		RELH1_5M:standard_name = "relative_humidity" ;
		RELH1_5M:long_name = "calculated relative humidity at 1.5 meters" ;
		RELH1_5M:units = "percent" ;
		RELH1_5M:_FillValue = -9999.f ;
		RELH1_5M:observation_type = "calculated" ;
		RELH1_5M:coordinates = "TIME LATITUDE LONGITUDE" ;
	float RELH2_0M(TIME) ;
		RELH2_0M:standard_name = "relative_humidity" ;
		RELH2_0M:long_name = "calculated relative humidity at 2.0 meters" ;
		RELH2_0M:units = "percent" ;
		RELH2_0M:_FillValue = -9999.f ;
		RELH2_0M:observation_type = "calculated" ;
		RELH2_0M:coordinates = "TIME LATITUDE LONGITUDE" ;
	char history(h_num, h_string) ;
		history:long_name = "file history information" ;

// global attributes:
		:project = "Integrated Marine Observing System (IMOS)" ;
		:conventions = "IMOS version 1.3" ;
		:title = "Heat and radiative flux data from Tangaroa" ;
		:institution = "Australian Bureau of Meteorology" ;
		:date_created = "2015-02-06T04:22:08Z" ;
		:comment = "COARE Bulk Flux Algorithm version 3.0b (Fairall et al.,2003: J.Climate,16,571-591)" ;
		:source = "Ship observation" ;
		:references = "http://www.imos.org.au" ;
		:netcdf_version = "3.6.1" ;
		:platform_code = "ZMFR" ;
		:naming_authority = "IMOS" ;
		:cdm_data_type = "Trajectory" ;
		:geospatial_lat_min = -67.671f ;
		:geospatial_lat_max = -67.1225f ;
		:geospatial_lon_min = 164.15f ;
		:geospatial_lon_max = 165.124f ;
		:geospatial_vertical_min = 0.f ;
		:geospatial_vertical_max = 0.f ;
		:time_coverage_start = "2015-02-05T00:01:00Z" ;
		:time_coverage_end = "2015-02-05T23:57:00Z" ;
		:data_centre = "eMarine Information Infrastructure (eMII)" ;
		:data_center_email = "info@emii.org.au" ;
		:author = "Ruslan Verein" ;
		:author_email = "r.verein@bom.gov.au" ;
		:principal_investigator = "Eric Schulz" ;
		:citation = "Citation to be used in publications should follow \n",
			"the format: \'IMOS.[year-of-data-download],[Title],[Data access URL],accessed \n",
			"[date-of access]\'" ;
		:acknowledgement = "Any users of IMOS data are required to clearly acknowledge the source of the material in the format: \"Data was sourced from the Integrated Marine Observing System (IMOS) - IMOS is supported by the Australian Government through the National Collaborative Research Infrastructure Strategy (NCRIS) and the Super Science Initiative (SSI).\"" ;
		:distribution_statement = "Data may be re-used, provided that related metadata explaining the data has been reviewed by the user, and the data is appropriately acknowledged. Data, products and services from IMOS are provided \"as is\" without any warranty as to fitness for a particular purpose." ;
		:file_version = "Level 2 - Derived product" ;
		:file_version_quality_control = "All data in this file has been \n",
			"through the BOM quality control procedure (Reference Table F) and was classed Z \n",
			"(passes all tests)" ;
		:site = "RV TANGAROA" ;
		:IMO = "9011571" ;
		:zi = "600.0" ;
		:zi_comment = "atmospheric boundary layer depth used in \n",
			"calculations, m" ;
		:jcool = "1" ;
		:jcool_comment = "1 - cool skin calculated, 0 - measured by IR \n",
			"radiometer" ;
		:jwarm = "1" ;
		:jwarm_comment = "1 - warm layer calculated, 0 - measured by IR \n",
			"radiometer" ;
		:jwave = "0" ;
		:jwave_comment = "wave state option: 0 - Charnock (Smith, 1988), \n",
			"1 - Oost et al. (2001), 2 - Taylor and Yelland (2000)" ;
		:data_comment = "for complete list of instruments see corresponding file version 1 (FV01)" ;
		:Conventions = "CF-1.6,IMOS-1.3" ;
		:data_centre_email = "info@emii.org.au" ;
		:history = "Wed Nov  4 16:19:27 2015: ncks -a -d TIME,,,10 self_referencing.nc temp.nc" ;
		:NCO = "4.4.2" ;
data:

 TIME = 23776.0013888888, 23776.0847222223, 23776.1194444443, 
    23776.1541666668, 23776.2062499998, 23776.2652777778, 23776.3034722223, 
    23776.3520833333, 23776.3937499998, 23776.4423611113, 23776.4909722223, 
    23776.5430555558, 23776.5777777778, 23776.6194444443, 23776.6576388888, 
    23776.6993055558, 23776.7618055558, 23776.8138888888, 23776.8555555558, 
    23776.8972222223, 23776.9423611113, 23776.9874999998 ;

 LATITUDE = -67.1658, -67.15, -67.1441, -67.138, -67.1232, -67.1491, 
    -67.2412, -67.2781, -67.4248, -67.5203, -67.6414, -67.6572, -67.5759, 
    -67.4863, -67.3765, -67.2966, -67.2032, -67.2667, -67.3479, -67.4999, 
    -67.6213, -67.5793 ;

 LONGITUDE = 164.189, 164.15, 164.16, 164.167, 164.165, 164.341, 164.222, 
    164.527, 164.408, 164.505, 164.663, 164.908, 165.049, 165.046, 165.001, 
    164.881, 164.715, 164.831, 165.029, 165.039, 164.968, 164.679 ;

 PL_CMP = 274, 131.9, 152.3, 156.8, 337.1, 290.9, 32.2, 14.1, 35.2, 45.8, 
    307.6, 216.2, 219.8, 176.1, 134.1, 104.4, 302.2, 346.1, 36.2, 2.8, 35.9, 
    158.1 ;

 PL_CRS = 274.1, 162.5, 218.5, 197.8, 177.7, 286.3, 35.8, 10.6, 37.3, 44.1, 
    308, 216.3, 216.9, 178.2, 132.6, 105.3, 296.9, 347.8, 35.4, 1.5, 32.7, 
    160.4 ;

 PL_SPD = 5.5, 0.4, 0.3, 0.3, 0.2, 3.3, 4.4, 5.2, 5.4, 5.2, 2.9, 3.5, 3.9, 
    3.5, 4.2, 5, 2.4, 4.6, 5.1, 5.4, 4.9, 5 ;

 WDIR = 181.2, 227.2, 218.6, 224.4, 241.4, 234, 234.8, 225.6, 260.9, 287.5, 
    298.7, 295.8, 269.7, 335.6, 66.7, 83.4, 244.8, 152.6, 14.3, 40.3, 278.8, 
    333.4 ;

 WSPD = 5.7, 7.3, 7.7, 7.2, 8.7, 8.7, 8.5, 8.5, 6.8, 6.9, 8.1, 12.9, 4.1, 
    2.2, 3.6, 2.7, 11.9, 2.6, 1.9, 5.7, 19.1, 10.8 ;

 WIND_H = 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24 ;

 WIND_FLAG = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 ATMP = 992.5, 993.1, 993.1, 993.2, 993.2, 993.2, 993.2, 993.1, 993.7, 993.3, 
    992.7, 991.6, 991.1, 990.8, 990.8, 990.6, 990.5, 989.8, 989.3, 988.6, 
    987.7, 988.4 ;

 ATMP_H = 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 
    12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5 ;

 ATMP_FLAG = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 AIRT = -0.6, -2.1, -2.6, -2.7, -1.8, -2.3, -2.3, -2.5, -3.6, -3.6, -3.1, -3, 
    -2.5, -2.7, -2.8, -2.9, -3.8, -1.8, -1.1, -1, -2.7, -3 ;

 AIRT_H = 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 
    14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6 ;

 AIRT_FLAG = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 RELH = 72.2, 73, 69.2, 66.2, 64.6, 73.4, 72, 73.6, 77.4, 76.6, 71.2, 67, 
    67.4, 72, 72, 72, 78, 67.8, 67.2, 64.6, 67.4, 69.2 ;

 RELH_H = 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 
    14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6, 14.6 ;

 RELH_FLAG = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 TEMP = -1.317, -1.0647, -1.231, -1.2592, -1.2971, -1.1264, -1.283, -1.3007, 
    -0.9275, -0.8478, -0.9581, -1.1155, -1.0789, -1.3118, -1.2316, -1.2269, 
    -1.3771, -1.3319, -1.166, -1.2084, -0.9597, -0.9644 ;

 TEMP_H = 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3 ;

 TEMP_FLAG = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 RAIN_AMOUNT = 0.1, 0, 0.6, 0, 0, 0, 0, 0.4, 0, 0.4, 0.7, 0.1, 0.1, 0.3, 0.8, 
    0, 1.5, 0.3, 0, 0, 0, 0.7 ;

 RAIN_AMOUNT_H = 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 
    18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2 ;

 RAIN_AMOUNT_FLAG = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1 ;

 SW = 738.7, 676.4, 657.9, 289.8, 476, 327.6, 193.1, 21.4, 3.7, 0, 0, 0, 0, 
    0, 0, 20.8, 121.8, 298.2, 374.4, 462, 578.2, 659.2 ;

 SW_H = 15.3, 15.3, 15.3, 15.3, 15.3, 15.3, 15.3, 15.3, 15.3, 15.3, 15.3, 
    15.3, 15.3, 15.3, 15.3, 15.3, 15.3, 15.3, 15.3, 15.3, 15.3, 15.3 ;

 SW_FLAG = 2, 1, 2, 2, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1 ;

 LW = 232.3, 222.7, 223.6, 233.3, 212.9, 217.6, 220.9, 288.9, 290.1, 287.7, 
    286.8, 263.9, 214.3, 215, 232.7, 221.3, 208.1, 211.8, 211.8, 221.2, 
    209.8, 256.1 ;

 LW_H = 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 
    18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2, 18.2 ;

 LW_FLAG = 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3 ;

 HS = -5.530089, 7.79121, 11.91465, 11.99592, 2.776049, 10.85179, 8.744937, 
    11.6972, 25.33899, 26.46922, 22.39748, 29.36836, 6.754734, 3.558745, 
    7.214238, 5.971715, 35.74469, 0.1135716, -0.508918, -2.726293, 40.16847, 
    26.82658 ;

 HL = 10.58714, 26.52441, 32.84274, 33.80349, 35.0185, 31.41995, 30.72651, 
    30.93284, 31.55755, 33.12394, 38.3847, 61.43007, 20.80054, 10.77139, 
    17.14229, 13.84296, 46.11297, 9.932697, 2.347661, 19.35552, 91.07937, 
    50.71571 ;

 H_RAIN = 0.06743633, 0, 1.677527, 0, 0, 0, 0, 0.9905027, 0, 1.500753, 
    2.424883, 0.3434108, 0.2816341, 0.7227817, 2.181409, 0, 5.009088, 
    0.5562372, 0, 0, 0, 2.425655 ;

 TAU = 0.02760131, 0.07178884, 0.08242486, 0.07153736, 0.1027948, 0.1067381, 
    0.1005441, 0.101765, 0.06697644, 0.06923894, 0.09534737, 0.2803872, 
    0.0221936, 0.007007649, 0.01752345, 0.01038743, 0.2325931, 0.008012, 
    0.001466323, 0.03459444, 0.7562687, 0.1812678 ;

 SST = -1.419884, -1.186227, -1.355034, -1.388387, -1.414505, -1.244392, 
    -1.400371, -1.357696, -1.016958, -0.942644, -1.040836, -1.19726, 
    -1.330503, -1.679, -1.462597, -1.534446, -1.495481, -1.627062, -1.513471, 
    -1.253734, -1.04151, -1.057681 ;

 HEAT_NET = -618.4614, -519.9753, -493.67, -154.3292, -318.6216, -177.713, 
    -57.30094, 42.34422, 73.68118, 82.53188, 84.15852, 135.6944, 119.9733, 
    104.5381, 98.34297, 84.88882, 64.46061, -178.2144, -257.8586, -333.9059, 
    -317.0894, -492.3223 ;

 MASS_NET = -0.0003374318, 1.060977e-05, -0.002036863, 1.35214e-05, 
    1.40074e-05, 1.256798e-05, 1.229061e-05, -0.001354294, 1.262302e-05, 
    -0.001353417, -0.002376313, -0.0003170946, -0.0003333465, -0.001020691, 
    -0.002726476, 5.537184e-06, -0.005106555, -0.001021027, 9.390645e-07, 
    7.742208e-06, 3.643175e-05, -0.00237138 ;

 LW_NET = 74.55302, 84.90702, 83.28809, 73.73241, 93.40387, 89.5973, 
    85.70711, 19.93719, 20.28113, 22.93871, 23.37635, 44.89599, 92.41799, 
    90.20799, 73.98644, 84.73015, 97.70395, 93.53828, 94.1106, 86.05492, 
    98.06178, 53.0794 ;

 SW_NET = -698.0715, -639.198, -621.7155, -273.861, -449.82, -309.582, 
    -182.4795, -20.223, -3.4965, 0, 0, 0, 0, 0, 0, -19.656, -115.101, 
    -281.799, -353.808, -436.59, -546.399, -622.944 ;

 WSPD10M = 5.380276, 6.808802, 7.17861, 6.719315, 8.093864, 8.095823, 
    7.911747, 7.912724, 6.360563, 6.453012, 7.550324, 11.91105, 3.856134, 
    2.092327, 3.395417, 2.563416, 11.01064, 2.439866, 1.835768, 5.341228, 
    17.44209, 10.01518 ;

 AIRT1_5M = -0.5663623, -1.796389, -2.226796, -2.30641, -1.610711, -1.975929, 
    -2.007138, -2.156601, -2.897816, -2.882483, -2.550548, -2.561066, 
    -2.09435, -2.311597, -2.340398, -2.4175, -3.255424, -1.650296, 
    -0.9428698, -0.9228774, -2.318043, -2.512998 ;

 AIRT2_0M = -0.5451934, -1.814793, -2.253026, -2.334741, -1.616199, 
    -1.996948, -2.024592, -2.179793, -2.959428, -2.945794, -2.596327, 
    -2.596151, -2.122947, -2.338218, -2.374696, -2.454219, -3.302247, 
    -1.6511, -0.9344332, -0.9135451, -2.347356, -2.552903 ;

 RELH1_5M = 74.54707, 79.61785, 77.18143, 75.15481, 71.44819, 79.84705, 
    78.4722, 80.22392, 86.85897, 86.36209, 80.30585, 75.02024, 77.48436, 
    81.43396, 81.58681, 82.11543, 85.11476, 75.21161, 65.48044, 70.0271, 
    74.23325, 77.59737 ;

 RELH2_0M = 74.1069, 78.85734, 76.27061, 74.14147, 70.62613, 79.09727, 
    77.71671, 79.45721, 85.81678, 85.28632, 79.28026, 74.06905, 76.38535, 
    80.414, 80.54738, 81.0219, 84.2849, 74.37967, 65.0431, 69.28867, 
    73.39404, 76.62269 ;

 history =
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;
}
