
netcdf Lake_Superior_-_Forecast_Forcing_-_2D_-_Current_Year_best {
dimensions:
    nsigma = 8 ;
    nx = 4 ;
    ny = 4 ;
    time = 4 ;
variables:
    float at(time, ny, nx) ;
        at:units = "Celsius" ;
        at:long_name = "Air Temperature" ;
        at:missing_value = -99999.f ;
        at:standard_name = "air_temperature" ;
        at:coordinates = "time_run time lat lon " ;
    float cl(time, ny, nx) ;
        cl:units = "fraction" ;
        cl:long_name = "Cloud cover" ;
        cl:missing_value = -99999.f ;
        cl:standard_name = "cloud_cover" ;
        cl:coordinates = "time_run time lat lon " ;
    float dp(time, ny, nx) ;
        dp:units = "Celsius" ;
        dp:long_name = "Dew Point" ;
        dp:missing_value = -99999.f ;
        dp:standard_name = "dew_point" ;
        dp:coordinates = "time_run time lat lon " ;
    float air_u(time, ny, nx) ;
        air_u:units = "m/s" ;
        air_u:long_name = "Eastward Air Velocity" ;
        air_u:missing_value = -99999.f ;
        air_u:standard_name = "eastward_wind" ;
        air_u:coordinates = "time_run time lat lon " ;
    float air_v(time, ny, nx) ;
        air_v:units = "m/s" ;
        air_v:long_name = "Northward Air Velocity" ;
        air_v:missing_value = -99999.f ;
        air_v:standard_name = "northward_wind" ;
        air_v:coordinates = "time_run time lat lon " ;
    double time_offset(time) ;
        time_offset:long_name = "offset hour from start of run for coordinate = time" ;
        time_offset:standard_name = "forecast_period" ;
        time_offset:units = "hours since 2016-01-01T12:00:00Z" ;
        time_offset:missing_value = NaN ;
    float lon(ny, nx) ;
        lon:units = "degrees_east" ;
        lon:long_name = "Longitude" ;
        lon:standard_name = "longitude" ;
        lon:_CoordinateAxisType = "Lon" ;
    float lat(ny, nx) ;
        lat:units = "degrees_north" ;
        lat:long_name = "Latitude" ;
        lat:standard_name = "latitude" ;
        lat:_CoordinateAxisType = "Lat" ;
    float depth(ny, nx) ;
        depth:units = "meters" ;
        depth:long_name = "Bathymetry" ;
        depth:positive = "down" ;
        depth:standard_name = "depth" ;
        depth:coordinates = "lat lon " ;
        depth:_CoordinateAxisType = "Height" ;
        depth:_CoordinateZisPositive = "down" ;
    float sigma(nsigma) ;
        sigma:units = "1" ;
        sigma:long_name = "Sigma Stretched Vertical Coordinate at Nodes" ;
        sigma:axis = "Z" ;
        sigma:positive = "down" ;
        sigma:standard_name = "ocean_sigma_coordinate" ;
        sigma:formula_terms = "sigma: sigma eta: eta depth: depth" ;
        sigma:_CoordinateAxisType = "GeoZ" ;
        sigma:_CoordinateZisPositive = "down" ;
        sigma:_CoordinateTransformType = "Vertical" ;
        sigma:_CoordinateAxes = "sigma" ;
    double time(time) ;
        time:long_name = "Forecast time for ForecastModelRunCollection" ;
        time:standard_name = "time" ;
        time:units = "hours since 2016-01-01T12:00:00Z" ;
        time:missing_value = NaN ;
        time:_CoordinateAxisType = "Time" ;
    double time_run(time) ;
        time_run:long_name = "run times for coordinate = time" ;
        time_run:standard_name = "forecast_reference_time" ;
        time_run:units = "hours since 2016-01-01T12:00:00Z" ;
        time_run:missing_value = NaN ;
        time_run:_CoordinateAxisType = "RunTime" ;

// global attributes:
        :institution = "NOAA/GLERL" ;
        :title = "Great Lakes Coastal Forecasting System (GLCFS), FORECAST" ;
        :data_source = "NDFD" ;
        :comment1 = "Lake Superior 10 km bathymetric grid" ;
        :comment2 = "1-hourly input data starting at validtime" ;
        :comment3 = "Generated 2x per day following the 0,12 Z Forecast runs" ;
        :validtime = "01-JAN-2016 00:00 GMT" ;
        :validtime_DOY = "001, 2016 00:00 GMT" ;
        :author = "gregory.lang@noaa.gov" ;
        :references = "http://www.glerl.noaa.gov/res/glcfs/" ;
        :creation_date = "Mon Nov  7 01:06:02 2016 GMT" ;
        :disclaimer = "http://www.glerl.noaa.gov/home/notice.html" ;
        :_CoordSysBuilder = "ucar.nc2.dataset.conv.CF1Convention" ;
        :Conventions = "CF-1.6" ;
        :cdm_data_type = "GRID" ;
        :featureType = "GRID" ;
        :location = "Proto fmrc:Lake_Superior_-_Forecast_Forcing_-_2D_-_Current_Year" ;
        :history = "FMRC Best Dataset" ;
}
