netcdf 2d-static-grid {
dimensions:
    lat = 2;
    lon = 2;
variables:
    double lat(lat);
        lat:standard_name = "latitude";
        lat:units = "degrees_north";
    double lon(lon);
        lon:standard_name = "longitude";
        lon:units = "degrees_east";
    double T(lat, lon);
        T:standard_name = "sea_water_temperature";
        T:units = "deg_C";
}
