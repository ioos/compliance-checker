
netcdf OCOS {
dimensions:
	Nuser = 25 ;
	boundary = 4 ;
	eta_psi = 3 ;
	eta_rho = 4 ;
	eta_u = 4 ;
	eta_v = 3 ;
	ocean_time = 2 ;
	s_rho = 2 ;
	s_w = 3 ;
	tracer = 2 ;
	xi_psi = 3 ;
	xi_rho = 4 ;
	xi_u = 3 ;
	xi_v = 4 ;
variables:
	int ntimes ;
		ntimes:long_name = "number of long time-steps" ;
	int ndtfast ;
		ndtfast:long_name = "number of short time-steps" ;
	double dt ;
		dt:long_name = "size of long time-steps" ;
		dt:units = "second" ;
	double dtfast ;
		dtfast:long_name = "size of short time-steps" ;
		dtfast:units = "second" ;
	double dstart ;
		dstart:long_name = "time stamp assigned to model initilization" ;
		dstart:units = "days since 2005-01-01 00:00:00" ;
	int nHIS ;
		nHIS:long_name = "number of time-steps between history records" ;
	int ndefHIS ;
		ndefHIS:long_name = "number of time-steps between the creation of history files" ;
	int nRST ;
		nRST:long_name = "number of time-steps between restart records" ;
	int ntsAVG ;
		ntsAVG:long_name = "starting time-step for accumulation of time-averaged fields" ;
	int nAVG ;
		nAVG:long_name = "number of time-steps between time-averaged records" ;
	int ndefAVG ;
		ndefAVG:long_name = "number of time-steps between the creation of average files" ;
	double Falpha ;
		Falpha:long_name = "Power-law shape barotropic filter parameter" ;
	double Fbeta ;
		Fbeta:long_name = "Power-law shape barotropic filter parameter" ;
	double Fgamma ;
		Fgamma:long_name = "Power-law shape barotropic filter parameter" ;
	double nl_tnu2(tracer) ;
		nl_tnu2:long_name = "nonlinear model Laplacian mixing coefficient for tracers" ;
		nl_tnu2:units = "meter2 second-1" ;
	double nl_visc2 ;
		nl_visc2:long_name = "nonlinear model Laplacian mixing coefficient for momentum" ;
		nl_visc2:units = "meter2 second-1" ;
	double Akt_bak(tracer) ;
		Akt_bak:long_name = "background vertical mixing coefficient for tracers" ;
		Akt_bak:units = "meter2 second-1" ;
	double Akv_bak ;
		Akv_bak:long_name = "background vertical mixing coefficient for momentum" ;
		Akv_bak:units = "meter2 second-1" ;
	double Akk_bak ;
		Akk_bak:long_name = "background vertical mixing coefficient for turbulent energy" ;
		Akk_bak:units = "meter2 second-1" ;
	double Akp_bak ;
		Akp_bak:long_name = "background vertical mixing coefficient for length scale" ;
		Akp_bak:units = "meter2 second-1" ;
	double rdrg ;
		rdrg:long_name = "linear drag coefficient" ;
		rdrg:units = "meter second-1" ;
	double rdrg2 ;
		rdrg2:long_name = "quadratic drag coefficient" ;
	double Zob ;
		Zob:long_name = "bottom roughness" ;
		Zob:units = "meter" ;
	double Zos ;
		Zos:long_name = "surface roughness" ;
		Zos:units = "meter" ;
	double Znudg ;
		Znudg:long_name = "free-surface nudging/relaxation inverse time scale" ;
		Znudg:units = "day-1" ;
	double M2nudg ;
		M2nudg:long_name = "2D momentum nudging/relaxation inverse time scale" ;
		M2nudg:units = "day-1" ;
	double M3nudg ;
		M3nudg:long_name = "3D momentum nudging/relaxation inverse time scale" ;
		M3nudg:units = "day-1" ;
	double Tnudg(tracer) ;
		Tnudg:long_name = "Tracers nudging/relaxation inverse time scale" ;
		Tnudg:units = "day-1" ;
	double FSobc_in(boundary) ;
		FSobc_in:long_name = "free-surface inflow, nudging inverse time scale" ;
		FSobc_in:units = "second-1" ;
	double FSobc_out(boundary) ;
		FSobc_out:long_name = "free-surface outflow, nudging inverse time scale" ;
		FSobc_out:units = "second-1" ;
	double M2obc_in(boundary) ;
		M2obc_in:long_name = "2D momentum inflow, nudging inverse time scale" ;
		M2obc_in:units = "second-1" ;
	double M2obc_out(boundary) ;
		M2obc_out:long_name = "2D momentum outflow, nudging inverse time scale" ;
		M2obc_out:units = "second-1" ;
	double Tobc_in(boundary, tracer) ;
		Tobc_in:long_name = "tracers inflow, nudging inverse time scale" ;
		Tobc_in:units = "second-1" ;
	double Tobc_out(boundary, tracer) ;
		Tobc_out:long_name = "tracers outflow, nudging inverse time scale" ;
		Tobc_out:units = "second-1" ;
	double M3obc_in(boundary) ;
		M3obc_in:long_name = "3D momentum inflow, nudging inverse time scale" ;
		M3obc_in:units = "second-1" ;
	double M3obc_out(boundary) ;
		M3obc_out:long_name = "3D momentum outflow, nudging inverse time scale" ;
		M3obc_out:units = "second-1" ;
	double rho0 ;
		rho0:long_name = "mean density used in Boussinesq approximation" ;
		rho0:units = "kilogram meter-3" ;
	double gamma2 ;
		gamma2:long_name = "slipperiness parameter" ;
	int LtracerSrc(tracer) ;
		LtracerSrc:long_name = "tracer point sources and sink activation switch" ;
		LtracerSrc:flag_values = 0, 1 ;
		LtracerSrc:flag_meanings = ".FALSE. .TRUE." ;
	int spherical ;
		spherical:long_name = "grid type logical switch" ;
		spherical:flag_values = 0, 1 ;
		spherical:flag_meanings = "Cartesian spherical" ;
	double xl ;
		xl:long_name = "domain length in the XI-direction" ;
		xl:units = "meter" ;
	double el ;
		el:long_name = "domain length in the ETA-direction" ;
		el:units = "meter" ;
	int Vtransform ;
		Vtransform:long_name = "vertical terrain-following transformation equation" ;
	int Vstretching ;
		Vstretching:long_name = "vertical terrain-following stretching function" ;
	double theta_s ;
		theta_s:long_name = "S-coordinate surface control parameter" ;
	double theta_b ;
		theta_b:long_name = "S-coordinate bottom control parameter" ;
	double Tcline ;
		Tcline:long_name = "S-coordinate surface/bottom layer width" ;
		Tcline:units = "meter" ;
	double hc ;
		hc:long_name = "S-coordinate parameter, critical depth" ;
		hc:units = "meter" ;
	double s_rho(s_rho) ;
		s_rho:long_name = "S-coordinate at RHO-points" ;
		s_rho:valid_min = -1. ;
		s_rho:valid_max = 0. ;
		s_rho:positive = "up" ;
		s_rho:standard_name = "ocean_s_coordinate_g2" ;
		s_rho:formula_terms = "s: s_rho C: Cs_r eta: zeta depth: h depth_c: hc" ;
		s_rho:field = "s_rho, scalar" ;
	double s_w(s_w) ;
		s_w:long_name = "S-coordinate at W-points" ;
		s_w:valid_min = -1. ;
		s_w:valid_max = 0. ;
		s_w:positive = "up" ;
		s_w:standard_name = "ocean_s_coordinate_g2" ;
		s_w:formula_terms = "s: s_w C: Cs_w eta: zeta depth: h depth_c: hc" ;
		s_w:field = "s_w, scalar" ;
	double Cs_r(s_rho) ;
		Cs_r:long_name = "S-coordinate stretching curves at RHO-points" ;
		Cs_r:valid_min = -1. ;
		Cs_r:valid_max = 0. ;
		Cs_r:field = "Cs_r, scalar" ;
	double Cs_w(s_w) ;
		Cs_w:long_name = "S-coordinate stretching curves at W-points" ;
		Cs_w:valid_min = -1. ;
		Cs_w:valid_max = 0. ;
		Cs_w:field = "Cs_w, scalar" ;
	double user(Nuser) ;
		user:long_name = "user generic parameters" ;
		user:field = "user, scalar" ;
	double h(eta_rho, xi_rho) ;
		h:long_name = "bathymetry at RHO-points" ;
		h:units = "meter" ;
		h:coordinates = "lon_rho lat_rho" ;
		h:field = "bath, scalar" ;
	double f(eta_rho, xi_rho) ;
		f:long_name = "Coriolis parameter at RHO-points" ;
		f:units = "second-1" ;
		f:coordinates = "lon_rho lat_rho" ;
		f:field = "coriolis, scalar" ;
	double pm(eta_rho, xi_rho) ;
		pm:long_name = "curvilinear coordinate metric in XI" ;
		pm:units = "meter-1" ;
		pm:coordinates = "lon_rho lat_rho" ;
		pm:field = "pm, scalar" ;
	double pn(eta_rho, xi_rho) ;
		pn:long_name = "curvilinear coordinate metric in ETA" ;
		pn:units = "meter-1" ;
		pn:coordinates = "lon_rho lat_rho" ;
		pn:field = "pn, scalar" ;
	double lon_rho(eta_rho, xi_rho) ;
		lon_rho:long_name = "longitude of RHO-points" ;
		lon_rho:units = "degree_east" ;
		lon_rho:standard_name = "longitude" ;
		lon_rho:field = "lon_rho, scalar" ;
	double lat_rho(eta_rho, xi_rho) ;
		lat_rho:long_name = "latitude of RHO-points" ;
		lat_rho:units = "degree_north" ;
		lat_rho:standard_name = "latitude" ;
		lat_rho:field = "lat_rho, scalar" ;
	double lon_u(eta_u, xi_u) ;
		lon_u:long_name = "longitude of U-points" ;
		lon_u:units = "degree_east" ;
		lon_u:standard_name = "longitude" ;
		lon_u:field = "lon_u, scalar" ;
	double lat_u(eta_u, xi_u) ;
		lat_u:long_name = "latitude of U-points" ;
		lat_u:units = "degree_north" ;
		lat_u:standard_name = "latitude" ;
		lat_u:field = "lat_u, scalar" ;
	double lon_v(eta_v, xi_v) ;
		lon_v:long_name = "longitude of V-points" ;
		lon_v:units = "degree_east" ;
		lon_v:standard_name = "longitude" ;
		lon_v:field = "lon_v, scalar" ;
	double lat_v(eta_v, xi_v) ;
		lat_v:long_name = "latitude of V-points" ;
		lat_v:units = "degree_north" ;
		lat_v:standard_name = "latitude" ;
		lat_v:field = "lat_v, scalar" ;
	double lon_psi(eta_psi, xi_psi) ;
		lon_psi:long_name = "longitude of PSI-points" ;
		lon_psi:units = "degree_east" ;
		lon_psi:standard_name = "longitude" ;
		lon_psi:field = "lon_psi, scalar" ;
	double lat_psi(eta_psi, xi_psi) ;
		lat_psi:long_name = "latitude of PSI-points" ;
		lat_psi:units = "degree_north" ;
		lat_psi:standard_name = "latitude" ;
		lat_psi:field = "lat_psi, scalar" ;
	double angle(eta_rho, xi_rho) ;
		angle:long_name = "angle between XI-axis and EAST" ;
		angle:units = "radians" ;
		angle:coordinates = "lon_rho lat_rho" ;
		angle:field = "angle, scalar" ;
	double mask_rho(eta_rho, xi_rho) ;
		mask_rho:long_name = "mask on RHO-points" ;
		mask_rho:flag_values = 0., 1. ;
		mask_rho:flag_meanings = "land water" ;
		mask_rho:coordinates = "lon_rho lat_rho" ;
	double mask_u(eta_u, xi_u) ;
		mask_u:long_name = "mask on U-points" ;
		mask_u:flag_values = 0., 1. ;
		mask_u:flag_meanings = "land water" ;
		mask_u:coordinates = "lon_u lat_u" ;
	double mask_v(eta_v, xi_v) ;
		mask_v:long_name = "mask on V-points" ;
		mask_v:flag_values = 0., 1. ;
		mask_v:flag_meanings = "land water" ;
		mask_v:coordinates = "lon_v lat_v" ;
	double mask_psi(eta_psi, xi_psi) ;
		mask_psi:long_name = "mask on psi-points" ;
		mask_psi:flag_values = 0., 1. ;
		mask_psi:flag_meanings = "land water" ;
		mask_psi:coordinates = "lon_psi lat_psi" ;
	double ocean_time(ocean_time) ;
		ocean_time:long_name = "time since initialization" ;
		ocean_time:units = "seconds since 2005-01-01 00:00:00" ;
		ocean_time:calendar = "gregorian" ;
		ocean_time:field = "time, scalar, series" ;
		ocean_time:standard_name = "time" ;
	float zeta(ocean_time, eta_rho, xi_rho) ;
		zeta:long_name = "free-surface" ;
		zeta:units = "meter" ;
		zeta:time = "ocean_time" ;
		zeta:coordinates = "lon_rho lat_rho ocean_time" ;
		zeta:field = "free-surface, scalar, series" ;
		zeta:_FillValue = 1.e+37f ;
	float ubar(ocean_time, eta_u, xi_u) ;
		ubar:long_name = "vertically integrated u-momentum component" ;
		ubar:units = "meter second-1" ;
		ubar:time = "ocean_time" ;
		ubar:coordinates = "lon_u lat_u ocean_time" ;
		ubar:field = "ubar-velocity, scalar, series" ;
		ubar:_FillValue = 1.e+37f ;
	float vbar(ocean_time, eta_v, xi_v) ;
		vbar:long_name = "vertically integrated v-momentum component" ;
		vbar:units = "meter second-1" ;
		vbar:time = "ocean_time" ;
		vbar:coordinates = "lon_v lat_v ocean_time" ;
		vbar:field = "vbar-velocity, scalar, series" ;
		vbar:_FillValue = 1.e+37f ;
	float u(ocean_time, s_rho, eta_u, xi_u) ;
		u:long_name = "u-momentum component" ;
		u:units = "meter second-1" ;
		u:time = "ocean_time" ;
		u:coordinates = "lon_u lat_u s_rho ocean_time" ;
		u:field = "u-velocity, scalar, series" ;
		u:_FillValue = 1.e+37f ;
	float v(ocean_time, s_rho, eta_v, xi_v) ;
		v:long_name = "v-momentum component" ;
		v:units = "meter second-1" ;
		v:time = "ocean_time" ;
		v:coordinates = "lon_v lat_v s_rho ocean_time" ;
		v:field = "v-velocity, scalar, series" ;
		v:_FillValue = 1.e+37f ;
	float w(ocean_time, s_w, eta_rho, xi_rho) ;
		w:long_name = "vertical momentum component" ;
		w:units = "meter second-1" ;
		w:time = "ocean_time" ;
		w:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		w:field = "w-velocity, scalar, series" ;
		w:_FillValue = 1.e+37f ;
	float temp(ocean_time, s_rho, eta_rho, xi_rho) ;
		temp:long_name = "potential temperature" ;
		temp:units = "degree_Celsius" ;
		temp:time = "ocean_time" ;
		temp:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		temp:field = "temperature, scalar, series" ;
		temp:_FillValue = 1.e+37f ;
		temp:standard_name = "sea_water_potential_temperature" ;
	float salt(ocean_time, s_rho, eta_rho, xi_rho) ;
		salt:long_name = "salinity" ;
		salt:time = "ocean_time" ;
		salt:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		salt:field = "salinity, scalar, series" ;
		salt:_FillValue = 1.e+37f ;
		salt:standard_name = "sea_water_salinity" ;
		salt:units = "1" ;
	float AKv(ocean_time, s_w, eta_rho, xi_rho) ;
		AKv:long_name = "vertical viscosity coefficient" ;
		AKv:units = "meter2 second-1" ;
		AKv:time = "ocean_time" ;
		AKv:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		AKv:field = "AKv, scalar, series" ;
	float AKt(ocean_time, s_w, eta_rho, xi_rho) ;
		AKt:long_name = "temperature vertical diffusion coefficient" ;
		AKt:units = "meter2 second-1" ;
		AKt:time = "ocean_time" ;
		AKt:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		AKt:field = "AKt, scalar, series" ;
	float AKs(ocean_time, s_w, eta_rho, xi_rho) ;
		AKs:long_name = "salinity vertical diffusion coefficient" ;
		AKs:units = "meter2 second-1" ;
		AKs:time = "ocean_time" ;
		AKs:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		AKs:field = "AKs, scalar, series" ;
	float tke(ocean_time, s_w, eta_rho, xi_rho) ;
		tke:long_name = "turbulent kinetic energy" ;
		tke:units = "meter2 second-2" ;
		tke:time = "ocean_time" ;
		tke:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		tke:field = "tke, scalar, series" ;
	float shflux(ocean_time, eta_rho, xi_rho) ;
		shflux:long_name = "surface net heat flux" ;
		shflux:units = "watt meter-2" ;
		shflux:negative_value = "upward flux, cooling" ;
		shflux:positive_value = "downward flux, heating" ;
		shflux:time = "ocean_time" ;
		shflux:coordinates = "lon_rho lat_rho ocean_time" ;
		shflux:field = "surface heat flux, scalar, series" ;
		shflux:_FillValue = 1.e+37f ;
	float latent(ocean_time, eta_rho, xi_rho) ;
		latent:long_name = "net latent heat flux" ;
		latent:units = "watt meter-2" ;
		latent:negative_value = "upward flux, cooling" ;
		latent:positive_value = "downward flux, heating" ;
		latent:time = "ocean_time" ;
		latent:coordinates = "lon_rho lat_rho ocean_time" ;
		latent:field = "latent heat flux, scalar, series" ;
		latent:_FillValue = 1.e+37f ;
	float sensible(ocean_time, eta_rho, xi_rho) ;
		sensible:long_name = "net sensible heat flux" ;
		sensible:units = "watt meter-2" ;
		sensible:negative_value = "upward flux, cooling" ;
		sensible:positive_value = "downward flux, heating" ;
		sensible:time = "ocean_time" ;
		sensible:coordinates = "lon_rho lat_rho ocean_time" ;
		sensible:field = "sensible heat flux, scalar, series" ;
		sensible:_FillValue = 1.e+37f ;
	float lwrad(ocean_time, eta_rho, xi_rho) ;
		lwrad:long_name = "net longwave radiation flux" ;
		lwrad:units = "watt meter-2" ;
		lwrad:negative_value = "upward flux, cooling" ;
		lwrad:positive_value = "downward flux, heating" ;
		lwrad:time = "ocean_time" ;
		lwrad:coordinates = "lon_rho lat_rho ocean_time" ;
		lwrad:field = "longwave radiation, scalar, series" ;
		lwrad:_FillValue = 1.e+37f ;
	float swrad(ocean_time, eta_rho, xi_rho) ;
		swrad:long_name = "solar shortwave radiation flux" ;
		swrad:units = "watt meter-2" ;
		swrad:negative_value = "upward flux, cooling" ;
		swrad:positive_value = "downward flux, heating" ;
		swrad:time = "ocean_time" ;
		swrad:coordinates = "lon_rho lat_rho ocean_time" ;
		swrad:field = "shortwave radiation, scalar, series" ;
		swrad:_FillValue = 1.e+37f ;

// global attributes:
		:file = "ocean_his_4329.nc" ;
		:format = "netCDF-3 64bit offset file" ;
		:Conventions = "Unidata Dataset Discovery v1.0, CF-1.4" ;
		:type = "ROMS/TOMS history file" ;
		:title = "Regional Ocean Modeling System (ROMS): Oregon Coast" ;
		:rst_file = "ocean_rst.nc" ;
		:his_base = "ocean_his" ;
		:avg_file = "ocean_avg.nc" ;
		:grd_file = "/home/aruba/vol1/serofeev/OW/Prm/grd_ow2km_03_smooth04_lana.nc" ;
		:ini_file = "ocean_rst_y.nc" ;
		:frc_file_01 = "/home/aruba/vol1/serofeev/OW/Prm/frc_wind_var.nc" ;
		:frc_file_02 = "/home/aruba/vol1/serofeev/OW/Prm//frc_ow2km_Swrad.nc" ;
		:frc_file_03 = "/home/aruba/vol1/serofeev/OW/Prm/frc_ow2km_Tair.nc" ;
		:frc_file_04 = "/home/aruba/vol1/serofeev/OW/Prm/frc_ow2km_Pair.nc" ;
		:frc_file_05 = "/home/aruba/vol1/serofeev/OW/Prm/frc_ow2km_Qair.nc" ;
		:frc_file_06 = "/home/aruba/vol1/serofeev/OW/Prm/frc_ow2km_Cloud.nc" ;
		:frc_file_07 = "/home/aruba/vol1/serofeev/OW/Prm/ow2km_CR.nc" ;
		:frc_file_08 = "/home/aruba/vol1/serofeev/OW/Prm/rivers_2014-2016.nc" ;
		:frc_file_09 = "/home/aruba/vol1/serofeev/OW/Prm/ow2km_tide.nc" ;
		:bry_file = "/home/aruba/vol1/serofeev/OW/Prm/orw2km_bc_hycom.nc" ;
		:script_file = "ocean1.in" ;
		:NLM_LBC = "\n",
			"EDGE:  WEST   SOUTH  EAST   NORTH  \n",
			"zeta:  Cha    Cha    Clo    Cha    \n",
			"ubar:  Fla    Fla    Clo    Fla    \n",
			"vbar:  Fla    Fla    Clo    Fla    \n",
			"u:     RadNud RadNud Clo    RadNud \n",
			"v:     RadNud RadNud Clo    RadNud \n",
			"temp:  RadNud RadNud Clo    RadNud \n",
			"salt:  RadNud RadNud Clo    RadNud \n",
			"tke:   Gra    Gra    Clo    Gra" ;
		:svn_url = "https://www.myroms.org/svn/src/trunk" ;
		:svn_rev = "631M" ;
		:code_dir = "/home/aruba/vol1/serofeev/ROMS_3.6" ;
		:header_dir = "/home/aruba/vol1/serofeev/ROMS_3.6/ROMS/Include" ;
		:header_file = "ak_or.h" ;
		:os = "Linux" ;
		:cpu = "x86_64" ;
		:compiler_system = "pgi" ;
		:compiler_command = "/usr/local/pgi/linux86-64/2012/mpi/mpich/bin/mpif90" ;
		:compiler_flags = " -O3 -Mfree" ;
		:tiling = "002x008" ;
		:history = "ROMS/TOMS, Version 3.6, Sunday - November 6, 2016 -  6:36:25 AM" ;
		:ana_file = "ROMS/Functionals/ana_btflux.h, ROMS/Functionals/ana_hmixcoef.h, ROMS/Functionals/ana_nudgcoef.h, ROMS/Functionals/ana_rain.h, ROMS/Functionals/ana_stflux.h" ;
		:CPP_options = "AK_OR, ADD_FSOBC, ADD_M2OBC, ANA_BSFLUX, ANA_BTFLUX, ANA_RAIN, ANA_SSFLUX, ASSUMED_SHAPE, AVERAGES, BULK_FLUXES, CURVGRID, DJ_GRADPS, DOUBLE_PRECISION, LONGWAVE, MASKING, MIX_S_TS, MIX_S_UV, MPI, MY25_MIXING, NONLINEAR, NONLIN_EOS, N2S2_HORAVG, POWER_LAW, PROFILE, K_GSCHEME, RADIATION_2D, !RST_SINGLE, SALINITY, SOLAR_SOURCE, SOLVE3D, SPLINES, SPONGE, SSH_TIDES, TS_U3HADVECTION, TS_C4VADVECTION, TS_DIF2, TS_PSOURCE, UV_ADV, UV_COR, UV_U3HADVECTION, UV_C4VADVECTION, UV_QDRAG, UV_PSOURCE, UV_TIDES, UV_VIS2, VAR_RHO_2D" ;
		:id = "OCOS_latest_aggregation" ;
		:cdm_data_type = "Grid" ;
		:naming_authority = "org.nanoos" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0, CF-1.4" ;
		:summary = "Regional Ocean Modeling System (ROMS) 3-day, 4-hourly forecast for the Oregon coast at approximately 3-km resolution. While considerable effort has been made to implement all model components in a thorough, correct, and accurate manner, numerous sources of error are possible. As such, please use these data with the caution appropriate for any ocean related activity." ;
		:keywords = "Oceans; Ocean Temperature; Potential Temperature, Oceans; Salinity/Density; Salinity, Oceans; Sea Surface Topography; Sea Surface Height, Oceans; sea_water_potential_temperature ;sea_water_temperature; sea_water_salinity; Ocean Circulation; Ocean Currents; x_sea_water_velocity; y_sea_water_velocity" ;
		:keywords_vocabulary = "GCMD Science Keywords" ;
		:standard_name_vocabulary = "CF-1.4" ;
		:comment = "Model runs produced by Dr. Alex Kurapov (kurapov@coas.oregonstate.edu)." ;
		:creator_email = "kurapov@coas.oregonstate.edu" ;
		:creator_name = "Alex Kurapov" ;
		:creator_url = "http://ceoas.oregonstate.edu/profile/kurapov/" ;
		:institution = "Oregon State University" ;
		:project = "Northwest Association of Networked Ocean Observing Systems (NANOOS) (http://nanoos.org)" ;
		:contributor_name = "Svetlana Erofeeva" ;
		:contributor_role = "distributor" ;
		:publisher_email = "serofeev@coas.oregonstate.edu" ;
		:publisher_name = "Northwest Association of Networked Ocean Observing Systems (NANOOS) " ;
		:publisher_url = "http://nanoos.org" ;
		:license = "The data may be used and redistributed for free but is not intended for legal use, since it may contain inaccuracies. Neither the data Contributor, Oregon State University, NANOOS, NOAA, State of Oregon nor the United States Government, nor any of their employees or contractors, makes any warranty, express or implied, including warranties of merchantability and fitness for a particular purpose, or assumes any legal liability for the accuracy, completeness, or usefulness, of this information." ;
		:acknowledgment = "Northwest Association of Networked Ocean Observing Systems (NANOOS) receives funding from the National Oceanic and Atmospheric Administration (NOAA) as a Regional Association within the U.S. Integrated Ocean Observing System (IOOS). " ;
		:source = "Regional Ocean Modeling System (ROMS), http://myroms.org" ;
		:references = "http://myroms.org, http://nanoos.org" ;
}
