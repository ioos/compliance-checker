netcdf chap2 {
dimensions:
    time = 16;
variables:
    ushort bad_dtype; // ushort or uint16 is an illegal type
    float bad\ name; // PLEASE DON'T DO THIS
    double not_unique;
    double NOT_UNIQUE;

    double temperature(time);
        temperature:_FillValue = -20.;
        temperature:valid_range = 0., 20.;
        temperature:units = "deg_C";

    float no_reason(time, time);

    double wind_speed(time);
        wind_speed:_FillValue = 12.;
        wind_speed:valid_min = 0.;
        wind_speed:valid_max = 20.;
        wind_speed:units = "knots";
    
    :title = "A succint description of what is in the dataset";
    :institution = "CF";
    :history = "history goes here";
    :Conventions = "ACDD-1.1, CF-1.6";
}
